VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO single_port_ram
  CLASS BLOCK ;
  FOREIGN single_port_ram ;
  ORIGIN 0.000 0.000 ;
  SIZE 236.380 BY 247.100 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 234.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 234.160 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 230.700 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 230.700 184.810 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 234.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 234.160 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 230.700 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 230.700 181.510 ;
    END
  END VPWR
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 112.790 243.100 113.070 247.100 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 128.890 243.100 129.170 247.100 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 232.380 119.040 236.380 119.640 ;
    END
  END addr[5]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END clk
  PIN data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 138.550 243.100 138.830 247.100 ;
    END
  END data[0]
  PIN data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 141.770 243.100 142.050 247.100 ;
    END
  END data[1]
  PIN data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END data[2]
  PIN data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END data[3]
  PIN data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END data[4]
  PIN data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END data[5]
  PIN data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END data[6]
  PIN data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 232.380 95.240 236.380 95.840 ;
    END
  END data[7]
  PIN q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 232.380 146.240 236.380 146.840 ;
    END
  END q[0]
  PIN q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 232.380 125.840 236.380 126.440 ;
    END
  END q[1]
  PIN q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 232.380 142.840 236.380 143.440 ;
    END
  END q[2]
  PIN q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 232.380 139.440 236.380 140.040 ;
    END
  END q[3]
  PIN q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 232.380 136.040 236.380 136.640 ;
    END
  END q[4]
  PIN q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 232.380 122.440 236.380 123.040 ;
    END
  END q[5]
  PIN q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 232.380 129.240 236.380 129.840 ;
    END
  END q[6]
  PIN q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 232.380 132.640 236.380 133.240 ;
    END
  END q[7]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 232.380 115.640 236.380 116.240 ;
    END
  END we
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 230.460 234.005 ;
      LAYER met1 ;
        RECT 5.520 10.640 230.850 234.160 ;
      LAYER met2 ;
        RECT 7.000 242.820 112.510 243.100 ;
        RECT 113.350 242.820 128.610 243.100 ;
        RECT 129.450 242.820 138.270 243.100 ;
        RECT 139.110 242.820 141.490 243.100 ;
        RECT 142.330 242.820 230.830 243.100 ;
        RECT 7.000 4.280 230.830 242.820 ;
        RECT 7.000 4.000 73.870 4.280 ;
        RECT 74.710 4.000 80.310 4.280 ;
        RECT 81.150 4.000 86.750 4.280 ;
        RECT 87.590 4.000 99.630 4.280 ;
        RECT 100.470 4.000 106.070 4.280 ;
        RECT 106.910 4.000 109.290 4.280 ;
        RECT 110.130 4.000 112.510 4.280 ;
        RECT 113.350 4.000 115.730 4.280 ;
        RECT 116.570 4.000 230.830 4.280 ;
      LAYER met3 ;
        RECT 4.000 228.840 232.380 234.085 ;
        RECT 4.400 227.440 232.380 228.840 ;
        RECT 4.000 147.240 232.380 227.440 ;
        RECT 4.000 145.840 231.980 147.240 ;
        RECT 4.000 143.840 232.380 145.840 ;
        RECT 4.000 142.440 231.980 143.840 ;
        RECT 4.000 140.440 232.380 142.440 ;
        RECT 4.000 139.040 231.980 140.440 ;
        RECT 4.000 137.040 232.380 139.040 ;
        RECT 4.000 135.640 231.980 137.040 ;
        RECT 4.000 133.640 232.380 135.640 ;
        RECT 4.000 132.240 231.980 133.640 ;
        RECT 4.000 130.240 232.380 132.240 ;
        RECT 4.000 128.840 231.980 130.240 ;
        RECT 4.000 126.840 232.380 128.840 ;
        RECT 4.000 125.440 231.980 126.840 ;
        RECT 4.000 123.440 232.380 125.440 ;
        RECT 4.000 122.040 231.980 123.440 ;
        RECT 4.000 120.040 232.380 122.040 ;
        RECT 4.000 118.640 231.980 120.040 ;
        RECT 4.000 116.640 232.380 118.640 ;
        RECT 4.000 115.240 231.980 116.640 ;
        RECT 4.000 96.240 232.380 115.240 ;
        RECT 4.000 94.840 231.980 96.240 ;
        RECT 4.000 10.715 232.380 94.840 ;
      LAYER met4 ;
        RECT 58.255 13.095 174.240 212.665 ;
        RECT 176.640 13.095 177.540 212.665 ;
        RECT 179.940 13.095 203.025 212.665 ;
  END
END single_port_ram
END LIBRARY

