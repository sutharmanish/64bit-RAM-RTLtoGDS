* NGSPICE file created from single_port_ram.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

.subckt single_port_ram VGND VPWR addr[0] addr[1] addr[2] addr[3] addr[4] addr[5]
+ clk data[0] data[1] data[2] data[3] data[4] data[5] data[6] data[7] q[0] q[1] q[2]
+ q[3] q[4] q[5] q[6] q[7] we
X_3155_ _1567_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__clkbuf_1
X_2106_ ram\[62\]\[5\] ram\[63\]\[5\] _0604_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__mux2_1
X_3086_ net267 _1327_ _1519_ VGND VGND VPWR VPWR _1527_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2037_ _0830_ _0831_ _0832_ _0606_ _0573_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_37_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2939_ _1404_ net83 _1442_ VGND VGND VPWR VPWR _1447_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold340 ram\[7\]\[2\] VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold351 ram\[19\]\[1\] VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 addr_reg\[1\] VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 ram\[62\]\[2\] VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 ram\[29\]\[5\] VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 ram\[63\]\[7\] VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Left_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3911_ clknet_leaf_25_clk _0011_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3842_ clknet_leaf_29_clk _0404_ VGND VGND VPWR VPWR ram\[55\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3773_ clknet_leaf_20_clk _0335_ VGND VGND VPWR VPWR ram\[46\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2724_ net163 _1325_ _1313_ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__mux2_1
X_2655_ _1286_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__clkbuf_1
X_2586_ _1249_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__clkbuf_1
X_3207_ net68 _1319_ _1592_ VGND VGND VPWR VPWR _1596_ sky130_fd_sc_hd__mux2_1
X_3138_ _1558_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3069_ net38 _1327_ _1510_ VGND VGND VPWR VPWR _1518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold170 ram\[59\]\[4\] VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 ram\[6\]\[2\] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 ram\[25\]\[6\] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2440_ _1165_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__clkbuf_1
X_2371_ _1123_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_39_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3825_ clknet_leaf_22_clk _0387_ VGND VGND VPWR VPWR ram\[52\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3756_ clknet_leaf_20_clk _0318_ VGND VGND VPWR VPWR ram\[44\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2707_ _1314_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3687_ clknet_leaf_12_clk _0249_ VGND VGND VPWR VPWR ram\[35\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2638_ _1277_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2569_ _1240_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_81_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1940_ _0602_ ram\[61\]\[2\] _0570_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1871_ ram\[32\]\[1\] ram\[33\]\[1\] ram\[34\]\[1\] ram\[35\]\[1\] _0576_ _0577_
+ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__mux4_1
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3610_ clknet_leaf_1_clk _0172_ VGND VGND VPWR VPWR ram\[26\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_3541_ clknet_leaf_41_clk _0103_ VGND VGND VPWR VPWR ram\[17\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3472_ clknet_leaf_13_clk _0034_ VGND VGND VPWR VPWR ram\[8\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2423_ _1081_ net288 _1150_ VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__mux2_1
X_2354_ _1051_ _1113_ VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__or2_4
X_2285_ _1069_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3808_ clknet_leaf_23_clk _0370_ VGND VGND VPWR VPWR ram\[50\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3739_ clknet_leaf_19_clk _0301_ VGND VGND VPWR VPWR ram\[42\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2070_ _0593_ ram\[8\]\[4\] VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__and2b_1
X_2972_ _1402_ net359 _1461_ VGND VGND VPWR VPWR _1465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1923_ _0602_ ram\[37\]\[2\] _0570_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1854_ _0555_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_12_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1785_ _0544_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3524_ clknet_leaf_9_clk _0086_ VGND VGND VPWR VPWR ram\[15\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3455_ clknet_leaf_39_clk _0017_ VGND VGND VPWR VPWR ram\[7\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2406_ net386 _1064_ _1139_ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__mux2_1
X_3386_ _1690_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__clkbuf_1
X_2337_ net137 _1048_ _1104_ VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2268_ net9 VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__buf_4
X_2199_ _0551_ _0991_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold41 ram\[16\]\[2\] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 ram\[62\]\[1\] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 ram\[56\]\[5\] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 ram\[28\]\[4\] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 ram\[32\]\[4\] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 ram\[56\]\[7\] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 ram\[29\]\[4\] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_18_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_5 _1315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3240_ _1613_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__clkbuf_1
X_3171_ _1544_ net432 _1572_ VGND VGND VPWR VPWR _1576_ sky130_fd_sc_hd__mux2_1
X_2122_ ram\[24\]\[5\] ram\[25\]\[5\] ram\[26\]\[5\] ram\[27\]\[5\] _0561_ _0634_
+ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__mux4_1
X_2053_ ram\[56\]\[4\] ram\[57\]\[4\] ram\[58\]\[4\] ram\[59\]\[4\] _0615_ _0553_
+ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_52_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2955_ _1402_ net456 _1452_ VGND VGND VPWR VPWR _1456_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1906_ _0702_ _0703_ _0704_ _0644_ _0563_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__o221a_1
X_2886_ _1417_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1837_ _0545_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__clkbuf_4
Xhold500 ram\[44\]\[2\] VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__dlygate4sd3_1
X_1768_ _0567_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__clkbuf_4
X_3507_ clknet_leaf_9_clk _0069_ VGND VGND VPWR VPWR ram\[13\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_3438_ _0530_ net463 _0531_ VGND VGND VPWR VPWR _1718_ sky130_fd_sc_hd__mux2_1
X_3369_ _1681_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_68_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput20 net20 VGND VGND VPWR VPWR q[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2740_ _1083_ net393 _1329_ VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__mux2_1
X_2671_ _1070_ net466 _1294_ VGND VGND VPWR VPWR _1295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3223_ _1604_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__clkbuf_1
X_3154_ _1544_ net398 _1563_ VGND VGND VPWR VPWR _1567_ sky130_fd_sc_hd__mux2_1
X_2105_ _0590_ ram\[61\]\[5\] _0591_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3085_ _1526_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__clkbuf_1
X_2036_ ram\[38\]\[4\] ram\[39\]\[4\] _0649_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2938_ _1446_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2869_ _1407_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold341 ram\[63\]\[4\] VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold330 ram\[2\]\[4\] VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold352 ram\[13\]\[5\] VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold385 ram\[56\]\[1\] VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 ram\[59\]\[1\] VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 ram\[14\]\[0\] VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 ram\[12\]\[5\] VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3910_ clknet_leaf_14_clk _0010_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3841_ clknet_leaf_22_clk _0403_ VGND VGND VPWR VPWR ram\[54\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3772_ clknet_leaf_20_clk _0334_ VGND VGND VPWR VPWR ram\[46\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2723_ net13 VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2654_ net184 _1181_ _1285_ VGND VGND VPWR VPWR _1286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2585_ _1070_ net121 _1248_ VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__mux2_1
X_3206_ _1595_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3137_ _1544_ net491 _1554_ VGND VGND VPWR VPWR _1558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3068_ _1517_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__clkbuf_1
X_2019_ _0573_ _0811_ _0815_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold171 ram\[54\]\[0\] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold160 ram\[36\]\[0\] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 ram\[7\]\[0\] VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 ram\[21\]\[0\] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2370_ net178 _1068_ _1115_ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3824_ clknet_leaf_23_clk _0386_ VGND VGND VPWR VPWR ram\[52\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3755_ clknet_leaf_20_clk _0317_ VGND VGND VPWR VPWR ram\[44\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2706_ net218 _1312_ _1313_ VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3686_ clknet_leaf_11_clk _0248_ VGND VGND VPWR VPWR ram\[35\]\[4\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2637_ net376 _1181_ _1276_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2568_ _1070_ net216 _1239_ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__mux2_1
X_2499_ net141 _1181_ _1202_ VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_Left_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Left_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1870_ _0666_ _0667_ _0668_ _0560_ _0573_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__o221a_1
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3540_ clknet_leaf_42_clk _0102_ VGND VGND VPWR VPWR ram\[17\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3471_ clknet_leaf_5_clk _0033_ VGND VGND VPWR VPWR ram\[8\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2422_ _1154_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__clkbuf_1
X_2353_ _0530_ _0535_ _0533_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__or3b_4
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2284_ net312 _1068_ _1054_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3807_ clknet_leaf_23_clk _0369_ VGND VGND VPWR VPWR ram\[50\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_1999_ _0596_ _0795_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__and2_1
X_3738_ clknet_leaf_19_clk _0300_ VGND VGND VPWR VPWR ram\[42\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3669_ clknet_leaf_11_clk _0231_ VGND VGND VPWR VPWR ram\[33\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2971_ _1464_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1922_ _0568_ ram\[36\]\[2\] VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__and2b_1
X_1853_ _0651_ ram\[25\]\[0\] _0652_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1784_ _0583_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3523_ clknet_leaf_9_clk _0085_ VGND VGND VPWR VPWR ram\[15\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_3454_ clknet_leaf_40_clk _0016_ VGND VGND VPWR VPWR ram\[7\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2405_ _1144_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_4_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3385_ _1068_ net342 _1682_ VGND VGND VPWR VPWR _1690_ sky130_fd_sc_hd__mux2_1
X_2336_ _1053_ _1092_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__nor2_4
X_2267_ _1057_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2198_ ram\[28\]\[7\] ram\[29\]\[7\] _0654_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold20 ram\[16\]\[7\] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 ram\[13\]\[1\] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 ram\[63\]\[0\] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 ram\[0\]\[3\] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 ram\[48\]\[5\] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 ram\[2\]\[1\] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 ram\[19\]\[7\] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 ram\[14\]\[2\] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_6 _1315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3170_ _1575_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__clkbuf_1
X_2121_ _0559_ _0915_ _0544_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__o21a_1
X_2052_ _0845_ _0846_ _0847_ _0606_ _0585_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2954_ _1455_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2885_ _1404_ net291 _1412_ VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__mux2_1
X_1905_ ram\[10\]\[1\] ram\[11\]\[1\] _0576_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1836_ _0631_ _0633_ _0635_ _0626_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__a22o_1
X_1767_ _0000_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__buf_4
Xhold501 ram\[51\]\[7\] VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__dlygate4sd3_1
X_3506_ clknet_leaf_8_clk _0068_ VGND VGND VPWR VPWR ram\[13\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3437_ _1717_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__clkbuf_1
X_3368_ _1068_ net396 _1673_ VGND VGND VPWR VPWR _1681_ sky130_fd_sc_hd__mux2_1
X_2319_ _1091_ _1094_ VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__nor2_4
X_3299_ _1644_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_68_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput21 net21 VGND VGND VPWR VPWR q[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2670_ _0535_ _1266_ _0530_ _0533_ VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__or4bb_4
X_3222_ _1542_ net240 _1601_ VGND VGND VPWR VPWR _1604_ sky130_fd_sc_hd__mux2_1
X_3153_ _1566_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2104_ _0600_ ram\[60\]\[5\] VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__and2b_1
XFILLER_0_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3084_ net279 _1325_ _1519_ VGND VGND VPWR VPWR _1526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2035_ _0602_ ram\[37\]\[4\] _0570_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2937_ _1402_ net26 _1442_ VGND VGND VPWR VPWR _1446_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2868_ _1406_ net271 _1396_ VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__mux2_1
X_1819_ _0555_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__buf_4
X_2799_ _1114_ _1348_ VGND VGND VPWR VPWR _1367_ sky130_fd_sc_hd__nor2_4
Xhold320 ram\[13\]\[6\] VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold342 ram\[25\]\[2\] VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 ram\[25\]\[0\] VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 ram\[42\]\[0\] VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 ram\[53\]\[3\] VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 ram\[28\]\[5\] VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold364 ram\[12\]\[4\] VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 ram\[5\]\[7\] VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3840_ clknet_leaf_29_clk _0402_ VGND VGND VPWR VPWR ram\[54\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_70_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3771_ clknet_leaf_19_clk _0333_ VGND VGND VPWR VPWR ram\[46\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2722_ _1324_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2653_ _1266_ _1113_ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__nor2_4
X_2584_ _1161_ _1238_ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__nand2_4
XFILLER_0_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3205_ net30 _1317_ _1592_ VGND VGND VPWR VPWR _1595_ sky130_fd_sc_hd__mux2_1
X_3136_ _1557_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__clkbuf_1
X_3067_ net61 _1325_ _1510_ VGND VGND VPWR VPWR _1517_ sky130_fd_sc_hd__mux2_1
X_2018_ _0812_ _0813_ _0814_ _0618_ _0563_ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__o221a_1
X_3969_ clknet_leaf_37_clk _0525_ VGND VGND VPWR VPWR addr_reg\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold150 ram\[57\]\[5\] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 ram\[26\]\[0\] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 ram\[16\]\[4\] VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 ram\[11\]\[7\] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 ram\[9\]\[4\] VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3823_ clknet_leaf_30_clk _0385_ VGND VGND VPWR VPWR ram\[52\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3754_ clknet_leaf_20_clk _0316_ VGND VGND VPWR VPWR ram\[44\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2705_ _1053_ _1113_ VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__nor2_4
XFILLER_0_42_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3685_ clknet_leaf_11_clk _0247_ VGND VGND VPWR VPWR ram\[35\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2636_ _1266_ _1200_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__nor2_4
XFILLER_0_2_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2567_ _1149_ _1238_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__nand2_4
XFILLER_0_57_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2498_ _1183_ _1201_ VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__nor2_4
XFILLER_0_4_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3119_ _1546_ net511 _1538_ VGND VGND VPWR VPWR _1547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3470_ clknet_leaf_10_clk _0032_ VGND VGND VPWR VPWR ram\[8\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2421_ _1079_ net457 _1150_ VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__mux2_1
X_2352_ _1112_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__clkbuf_1
X_2283_ net14 VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3806_ clknet_leaf_23_clk _0368_ VGND VGND VPWR VPWR ram\[50\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_1998_ ram\[56\]\[3\] ram\[57\]\[3\] ram\[58\]\[3\] ram\[59\]\[3\] _0615_ _0553_
+ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3737_ clknet_leaf_24_clk _0299_ VGND VGND VPWR VPWR ram\[41\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3668_ clknet_leaf_11_clk _0230_ VGND VGND VPWR VPWR ram\[33\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3599_ clknet_leaf_1_clk _0161_ VGND VGND VPWR VPWR ram\[24\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2619_ _1266_ _1092_ VGND VGND VPWR VPWR _1267_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_7_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2970_ _1400_ net446 _1461_ VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__mux2_1
X_1921_ _0546_ _0714_ _0716_ _0718_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__a22o_1
X_1852_ _0549_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__buf_4
XFILLER_0_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1783_ _0004_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3522_ clknet_leaf_8_clk _0084_ VGND VGND VPWR VPWR ram\[15\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3453_ clknet_leaf_40_clk _0015_ VGND VGND VPWR VPWR ram\[7\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2404_ net387 _1062_ _1139_ VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__mux2_1
X_3384_ _1689_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_4_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2335_ _1103_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__clkbuf_1
X_2266_ net160 _1056_ _1054_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__mux2_1
X_2197_ _0659_ _0947_ _0961_ _0975_ _0990_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__a32o_1
XFILLER_0_62_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold21 ram\[6\]\[1\] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 ram\[39\]\[6\] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 ram\[33\]\[5\] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 ram\[3\]\[0\] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 ram\[20\]\[0\] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 ram\[28\]\[3\] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 ram\[16\]\[3\] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 ram\[22\]\[0\] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 ram\[41\]\[6\] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_7 _1317_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2120_ ram\[30\]\[5\] ram\[31\]\[5\] _0608_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__mux2_1
X_2051_ ram\[62\]\[4\] ram\[63\]\[4\] _0604_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2953_ _1400_ net273 _1452_ VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1904_ _0641_ ram\[9\]\[1\] _0550_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_60_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2884_ _1416_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__clkbuf_1
X_1835_ ram\[16\]\[0\] ram\[17\]\[0\] ram\[18\]\[0\] ram\[19\]\[0\] _0588_ _0634_
+ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__mux4_2
Xhold502 ram\[17\]\[5\] VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1766_ _0546_ _0552_ _0558_ _0565_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__a22o_1
X_3505_ clknet_leaf_13_clk _0067_ VGND VGND VPWR VPWR ram\[12\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3436_ net332 net14 _1709_ VGND VGND VPWR VPWR _1717_ sky130_fd_sc_hd__mux2_1
X_3367_ _1680_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__clkbuf_1
X_2318_ _1093_ VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__clkbuf_8
X_3298_ _1550_ net255 _1637_ VGND VGND VPWR VPWR _1644_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2249_ ram\[38\]\[7\] ram\[39\]\[7\] _0733_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput22 net22 VGND VGND VPWR VPWR q[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3221_ _1603_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__clkbuf_1
X_3152_ _1542_ net85 _1563_ VGND VGND VPWR VPWR _1566_ sky130_fd_sc_hd__mux2_1
X_2103_ _0893_ _0897_ _0003_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__o21ba_1
X_3083_ _1525_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__clkbuf_1
X_2034_ _0568_ ram\[36\]\[4\] VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2936_ _1445_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2867_ net12 VGND VGND VPWR VPWR _1406_ sky130_fd_sc_hd__buf_2
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1818_ _0559_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__clkbuf_4
Xhold310 ram\[42\]\[6\] VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__dlygate4sd3_1
X_2798_ _1366_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1749_ _0001_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__clkbuf_4
Xhold343 ram\[63\]\[6\] VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold332 ram\[31\]\[0\] VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 ram\[39\]\[2\] VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 ram\[19\]\[6\] VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 ram\[18\]\[1\] VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 ram\[31\]\[6\] VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 ram\[39\]\[1\] VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__dlygate4sd3_1
X_3419_ _1068_ net98 _1700_ VGND VGND VPWR VPWR _1708_ sky130_fd_sc_hd__mux2_1
Xhold398 ram\[14\]\[7\] VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3770_ clknet_leaf_20_clk _0332_ VGND VGND VPWR VPWR ram\[46\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2721_ net360 _1323_ _1313_ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2652_ _1284_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2583_ _1247_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__clkbuf_1
X_3204_ _1594_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__clkbuf_1
X_3135_ _1542_ net503 _1554_ VGND VGND VPWR VPWR _1557_ sky130_fd_sc_hd__mux2_1
X_3066_ _1516_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2017_ ram\[10\]\[3\] ram\[11\]\[3\] _0576_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__mux2_1
X_3968_ clknet_leaf_37_clk _0524_ VGND VGND VPWR VPWR addr_reg\[0\] sky130_fd_sc_hd__dfxtp_1
X_2919_ net196 _1319_ _1432_ VGND VGND VPWR VPWR _1436_ sky130_fd_sc_hd__mux2_1
X_3899_ clknet_leaf_33_clk _0461_ VGND VGND VPWR VPWR ram\[62\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold140 ram\[2\]\[6\] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 ram\[24\]\[4\] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 ram\[44\]\[7\] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 ram\[2\]\[0\] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 ram\[40\]\[5\] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 ram\[40\]\[3\] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3822_ clknet_leaf_31_clk _0384_ VGND VGND VPWR VPWR ram\[52\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3753_ clknet_leaf_21_clk _0315_ VGND VGND VPWR VPWR ram\[43\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2704_ net7 VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3684_ clknet_leaf_11_clk _0246_ VGND VGND VPWR VPWR ram\[35\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2635_ _1275_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2566_ _0537_ _1124_ _0540_ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__nor3_4
XFILLER_0_49_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2497_ _1051_ _1200_ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__or2_4
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3118_ net11 VGND VGND VPWR VPWR _1546_ sky130_fd_sc_hd__buf_2
X_3049_ _1506_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_81_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2420_ _1153_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__clkbuf_1
X_2351_ net237 _1068_ _1104_ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__mux2_1
X_2282_ _1067_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1997_ _0791_ _0792_ _0793_ _0606_ _0585_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__o221a_1
X_3805_ clknet_leaf_23_clk _0367_ VGND VGND VPWR VPWR ram\[50\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3736_ clknet_leaf_25_clk _0298_ VGND VGND VPWR VPWR ram\[41\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3667_ clknet_leaf_17_clk _0229_ VGND VGND VPWR VPWR ram\[33\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3598_ clknet_leaf_0_clk _0160_ VGND VGND VPWR VPWR ram\[24\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2618_ _1051_ _1089_ _1124_ _0540_ VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_7_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2549_ _1138_ _1183_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__nor2_4
XFILLER_0_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1920_ _0560_ _0717_ _0564_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__o21a_1
X_1851_ _0555_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3521_ clknet_leaf_13_clk _0083_ VGND VGND VPWR VPWR ram\[14\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_1782_ _0543_ _0566_ _0580_ _0581_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3452_ clknet_leaf_41_clk _0014_ VGND VGND VPWR VPWR ram\[7\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3383_ _1066_ net57 _1682_ VGND VGND VPWR VPWR _1689_ sky130_fd_sc_hd__mux2_1
X_2403_ _1143_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__clkbuf_1
X_2334_ net322 _1068_ _1095_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2265_ net8 VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__buf_4
X_2196_ _0581_ _0982_ _0989_ _0005_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__o31a_1
XFILLER_0_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3719_ clknet_leaf_41_clk _0281_ VGND VGND VPWR VPWR ram\[3\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold11 ram\[16\]\[6\] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 ram\[38\]\[6\] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 ram\[23\]\[2\] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 ram\[42\]\[7\] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 ram\[34\]\[5\] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 ram\[47\]\[6\] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 ram\[23\]\[3\] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 ram\[9\]\[5\] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 ram\[9\]\[0\] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_8 _1321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2050_ _0590_ ram\[61\]\[4\] _0591_ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_17_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2952_ _1454_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__clkbuf_1
X_1903_ _0604_ ram\[8\]\[1\] VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_60_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2883_ _1402_ net58 _1412_ VGND VGND VPWR VPWR _1416_ sky130_fd_sc_hd__mux2_1
X_1834_ _0549_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__buf_4
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1765_ _0560_ _0562_ _0564_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__o21a_1
X_3504_ clknet_leaf_13_clk _0066_ VGND VGND VPWR VPWR ram\[12\]\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold503 ram\[47\]\[3\] VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__dlygate4sd3_1
X_3435_ _1716_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3366_ _1066_ net366 _1673_ VGND VGND VPWR VPWR _1680_ sky130_fd_sc_hd__mux2_1
X_3297_ _1643_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__clkbuf_1
X_2317_ _1051_ _1092_ VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2248_ _0568_ ram\[37\]\[7\] _0577_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_68_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2179_ _0944_ _0972_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput23 net23 VGND VGND VPWR VPWR q[7] sky130_fd_sc_hd__buf_2
XFILLER_0_81_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3220_ _1540_ net467 _1601_ VGND VGND VPWR VPWR _1603_ sky130_fd_sc_hd__mux2_1
X_3151_ _1565_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2102_ _0894_ _0895_ _0896_ _0595_ _0596_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__o221a_1
X_3082_ net156 _1323_ _1519_ VGND VGND VPWR VPWR _1525_ sky130_fd_sc_hd__mux2_1
X_2033_ _0546_ _0824_ _0826_ _0828_ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2935_ _1400_ net304 _1442_ VGND VGND VPWR VPWR _1445_ sky130_fd_sc_hd__mux2_1
X_2866_ _1405_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__clkbuf_1
X_1817_ _0614_ _0616_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold300 ram\[48\]\[3\] VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 ram\[57\]\[7\] VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__dlygate4sd3_1
X_2797_ net239 _1327_ _1358_ VGND VGND VPWR VPWR _1366_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_15_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold333 ram\[51\]\[5\] VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 ram\[56\]\[6\] VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__dlygate4sd3_1
X_1748_ _0547_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__buf_4
Xhold322 ram\[31\]\[3\] VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 ram\[2\]\[7\] VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 ram\[49\]\[1\] VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 ram\[38\]\[7\] VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__dlygate4sd3_1
X_3418_ _1707_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__clkbuf_1
Xhold399 ram\[48\]\[2\] VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 ram\[62\]\[6\] VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3349_ net341 net13 _1664_ VGND VGND VPWR VPWR _1671_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2720_ net12 VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__buf_4
XFILLER_0_66_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2651_ net36 _1198_ _1276_ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2582_ _1087_ net101 _1239_ VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3203_ net408 _1315_ _1592_ VGND VGND VPWR VPWR _1594_ sky130_fd_sc_hd__mux2_1
X_3134_ _1556_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__clkbuf_1
X_3065_ net87 _1323_ _1510_ VGND VGND VPWR VPWR _1516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2016_ _0641_ ram\[9\]\[3\] _0550_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3967_ clknet_leaf_15_clk _0523_ VGND VGND VPWR VPWR ram\[39\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2918_ _1435_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3898_ clknet_leaf_32_clk _0460_ VGND VGND VPWR VPWR ram\[62\]\[0\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_30_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_45_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2849_ net213 _1327_ _1386_ VGND VGND VPWR VPWR _1394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold141 ram\[3\]\[6\] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 ram\[6\]\[0\] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold130 ram\[26\]\[4\] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 ram\[16\]\[5\] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 ram\[6\]\[7\] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 addr_reg\[3\] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 ram\[29\]\[3\] VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_21_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_54 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3821_ clknet_leaf_30_clk _0383_ VGND VGND VPWR VPWR ram\[52\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3752_ clknet_leaf_21_clk _0314_ VGND VGND VPWR VPWR ram\[43\]\[6\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_12_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_2
X_3683_ clknet_leaf_11_clk _0245_ VGND VGND VPWR VPWR ram\[35\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2703_ _1311_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2634_ net301 _1198_ _1267_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__mux2_1
X_2565_ _1237_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__clkbuf_1
X_2496_ _0533_ _0535_ _0530_ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__or3b_4
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3117_ _1545_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_38_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3048_ _1408_ net122 _1499_ VGND VGND VPWR VPWR _1506_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_438 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Left_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2350_ _1111_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__clkbuf_1
X_2281_ net327 _1066_ _1054_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_63_Left_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_1_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_72_Left_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1996_ ram\[62\]\[3\] ram\[63\]\[3\] _0604_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__mux2_1
X_3804_ clknet_leaf_23_clk _0366_ VGND VGND VPWR VPWR ram\[50\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3735_ clknet_leaf_24_clk _0297_ VGND VGND VPWR VPWR ram\[41\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3666_ clknet_leaf_11_clk _0228_ VGND VGND VPWR VPWR ram\[33\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3597_ clknet_leaf_44_clk _0159_ VGND VGND VPWR VPWR ram\[24\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2617_ _1265_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_81_Left_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2548_ _1228_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__clkbuf_1
X_2479_ net64 _1188_ _1184_ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1850_ _0649_ ram\[24\]\[0\] VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__and2b_1
XFILLER_0_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1781_ _0004_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3520_ clknet_leaf_4_clk _0082_ VGND VGND VPWR VPWR ram\[14\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3451_ clknet_leaf_39_clk _0013_ VGND VGND VPWR VPWR ram\[7\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3382_ _1688_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__clkbuf_1
X_2402_ net462 _1060_ _1139_ VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__mux2_1
X_2333_ _1102_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_4_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2264_ _1055_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2195_ _0986_ _0988_ _0003_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_7_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1979_ _0568_ ram\[36\]\[3\] VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__and2b_1
X_3718_ clknet_leaf_41_clk _0280_ VGND VGND VPWR VPWR ram\[3\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3649_ clknet_leaf_14_clk _0211_ VGND VGND VPWR VPWR ram\[30\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold12 ram\[57\]\[6\] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 ram\[49\]\[7\] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 ram\[58\]\[5\] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 ram\[56\]\[3\] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 ram\[59\]\[6\] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 ram\[17\]\[7\] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 ram\[21\]\[7\] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 ram\[36\]\[1\] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_54_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_9 _1323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2951_ _1398_ net395 _1452_ VGND VGND VPWR VPWR _1454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1902_ ram\[12\]\[1\] ram\[13\]\[1\] ram\[14\]\[1\] ram\[15\]\[1\] _0638_ _0624_
+ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2882_ _1415_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__clkbuf_1
X_1833_ _0618_ _0632_ _0544_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__o21a_1
X_1764_ _0563_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__clkbuf_4
Xhold504 ram\[19\]\[5\] VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3503_ clknet_leaf_8_clk _0065_ VGND VGND VPWR VPWR ram\[12\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3434_ net33 net13 _1709_ VGND VGND VPWR VPWR _1716_ sky130_fd_sc_hd__mux2_1
X_3365_ _1679_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3296_ _1548_ net515 _1637_ VGND VGND VPWR VPWR _1643_ sky130_fd_sc_hd__mux2_1
X_2316_ net1 net2 net3 VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__or3_4
X_2247_ _0561_ ram\[36\]\[7\] VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_68_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2178_ ram\[48\]\[6\] ram\[49\]\[6\] ram\[50\]\[6\] ram\[51\]\[6\] _0629_ _0652_
+ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3150_ _1540_ net361 _1563_ VGND VGND VPWR VPWR _1565_ sky130_fd_sc_hd__mux2_1
X_3081_ _1524_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__clkbuf_1
X_2101_ ram\[50\]\[5\] ram\[51\]\[5\] _0733_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__mux2_1
X_2032_ _0560_ _0827_ _0564_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2934_ _1444_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__clkbuf_1
X_2865_ _1404_ net477 _1396_ VGND VGND VPWR VPWR _1405_ sky130_fd_sc_hd__mux2_1
X_1816_ ram\[4\]\[0\] ram\[5\]\[0\] _0615_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2796_ _1365_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__clkbuf_1
Xhold301 ram\[43\]\[5\] VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__dlygate4sd3_1
X_1747_ _0000_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__buf_4
Xhold312 ram\[25\]\[1\] VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 ram\[23\]\[5\] VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 ram\[27\]\[1\] VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 ram\[60\]\[7\] VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 ram\[45\]\[7\] VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 ram\[8\]\[2\] VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 ram\[39\]\[0\] VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__dlygate4sd3_1
X_3417_ _1066_ net399 _1700_ VGND VGND VPWR VPWR _1707_ sky130_fd_sc_hd__mux2_1
Xhold389 ram\[3\]\[1\] VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__dlygate4sd3_1
X_3348_ _1670_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3279_ _1548_ net314 _1628_ VGND VGND VPWR VPWR _1634_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2650_ _1283_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2581_ _1246_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3202_ _1593_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_78_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3133_ _1540_ net254 _1554_ VGND VGND VPWR VPWR _1556_ sky130_fd_sc_hd__mux2_1
X_3064_ _1515_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2015_ _0593_ ram\[8\]\[3\] VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__and2b_1
XFILLER_0_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3966_ clknet_leaf_25_clk _0522_ VGND VGND VPWR VPWR ram\[39\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2917_ net299 _1317_ _1432_ VGND VGND VPWR VPWR _1435_ sky130_fd_sc_hd__mux2_1
X_3897_ clknet_leaf_28_clk _0459_ VGND VGND VPWR VPWR ram\[61\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2848_ _1393_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2779_ _1356_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold131 ram\[5\]\[1\] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 ram\[17\]\[1\] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 ram\[30\]\[2\] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 ram\[22\]\[4\] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 ram\[26\]\[5\] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 ram\[29\]\[1\] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 ram\[33\]\[3\] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 ram\[3\]\[7\] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3820_ clknet_leaf_30_clk _0382_ VGND VGND VPWR VPWR ram\[52\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3751_ clknet_leaf_21_clk _0313_ VGND VGND VPWR VPWR ram\[43\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_30_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2702_ net128 _1198_ _1303_ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3682_ clknet_leaf_11_clk _0244_ VGND VGND VPWR VPWR ram\[35\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2633_ _1274_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2564_ net169 _1198_ _1229_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2495_ _1199_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3116_ _1544_ net415 _1538_ VGND VGND VPWR VPWR _1545_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3047_ _1505_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3949_ clknet_leaf_27_clk _0505_ VGND VGND VPWR VPWR ram\[49\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2280_ net13 VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3803_ clknet_leaf_23_clk _0365_ VGND VGND VPWR VPWR ram\[50\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_1995_ _0602_ ram\[61\]\[3\] _0570_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3734_ clknet_leaf_18_clk _0296_ VGND VGND VPWR VPWR ram\[41\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3665_ clknet_leaf_15_clk _0227_ VGND VGND VPWR VPWR ram\[32\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2616_ net50 _1198_ _1257_ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3596_ clknet_leaf_44_clk _0158_ VGND VGND VPWR VPWR ram\[24\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2547_ net370 _1198_ _1220_ VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__mux2_1
X_2478_ net9 VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1780_ _0574_ _0579_ _0542_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_12_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3450_ clknet_leaf_39_clk _0012_ VGND VGND VPWR VPWR ram\[7\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_3381_ _1064_ net413 _1682_ VGND VGND VPWR VPWR _1688_ sky130_fd_sc_hd__mux2_1
X_2401_ _1142_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__clkbuf_1
X_2332_ net348 _1066_ _1095_ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2263_ net205 _1048_ _1054_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__mux2_1
X_2194_ _0944_ _0987_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_52 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3717_ clknet_leaf_40_clk _0279_ VGND VGND VPWR VPWR ram\[3\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_1978_ _0546_ _0770_ _0772_ _0774_ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3648_ clknet_leaf_3_clk _0210_ VGND VGND VPWR VPWR ram\[30\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3579_ clknet_leaf_2_clk _0141_ VGND VGND VPWR VPWR ram\[22\]\[1\] sky130_fd_sc_hd__dfxtp_1
Xhold13 ram\[25\]\[7\] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 ram\[55\]\[4\] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 ram\[38\]\[3\] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 ram\[41\]\[0\] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 ram\[57\]\[3\] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 ram\[28\]\[6\] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 ram\[28\]\[2\] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_54_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2950_ _1453_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__clkbuf_1
X_1901_ _0696_ _0698_ _0699_ _0626_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__a22o_1
X_2881_ _1400_ net142 _1412_ VGND VGND VPWR VPWR _1415_ sky130_fd_sc_hd__mux2_1
X_1832_ ram\[22\]\[0\] ram\[23\]\[0\] _0608_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1763_ _0002_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__clkinv_4
X_3502_ clknet_leaf_10_clk _0064_ VGND VGND VPWR VPWR ram\[12\]\[4\] sky130_fd_sc_hd__dfxtp_1
Xhold505 ram\[11\]\[2\] VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__dlygate4sd3_1
X_3433_ _1715_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__clkbuf_1
X_3364_ _1064_ net147 _1673_ VGND VGND VPWR VPWR _1679_ sky130_fd_sc_hd__mux2_1
X_3295_ _1642_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__clkbuf_1
X_2315_ _1090_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__buf_4
XFILLER_0_57_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2246_ _1034_ _1038_ _0542_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2177_ _0968_ _0969_ _0970_ _0595_ _0585_ VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__o221a_1
XFILLER_0_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3080_ net246 _1321_ _1519_ VGND VGND VPWR VPWR _1524_ sky130_fd_sc_hd__mux2_1
X_2100_ _0568_ ram\[49\]\[5\] _0591_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__a21o_1
X_2031_ ram\[42\]\[4\] ram\[43\]\[4\] _0651_ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2933_ _1398_ net340 _1442_ VGND VGND VPWR VPWR _1444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2864_ net11 VGND VGND VPWR VPWR _1404_ sky130_fd_sc_hd__buf_2
X_1815_ _0000_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__buf_4
X_2795_ net202 _1325_ _1358_ VGND VGND VPWR VPWR _1365_ sky130_fd_sc_hd__mux2_1
Xhold302 ram\[56\]\[0\] VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1746_ _0545_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__clkbuf_4
Xhold313 ram\[18\]\[2\] VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 ram\[25\]\[5\] VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold335 ram\[52\]\[6\] VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 ram\[27\]\[7\] VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 ram\[38\]\[5\] VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 ram\[15\]\[3\] VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__dlygate4sd3_1
X_3416_ _1706_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__clkbuf_1
Xhold379 ram\[46\]\[6\] VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__dlygate4sd3_1
X_3347_ net159 net12 _1664_ VGND VGND VPWR VPWR _1670_ sky130_fd_sc_hd__mux2_1
X_3278_ _1633_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_28_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2229_ ram\[58\]\[7\] ram\[59\]\[7\] _0556_ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2580_ _1085_ net115 _1239_ VGND VGND VPWR VPWR _1246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3201_ net325 _1312_ _1592_ VGND VGND VPWR VPWR _1593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3132_ _1555_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_78_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3063_ net272 _1321_ _1510_ VGND VGND VPWR VPWR _1515_ sky130_fd_sc_hd__mux2_1
X_2014_ ram\[12\]\[3\] ram\[13\]\[3\] ram\[14\]\[3\] ram\[15\]\[3\] _0600_ _0624_
+ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__mux4_1
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3965_ clknet_leaf_15_clk _0521_ VGND VGND VPWR VPWR ram\[39\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2916_ _1434_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3896_ clknet_leaf_28_clk _0458_ VGND VGND VPWR VPWR ram\[61\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2847_ net132 _1325_ _1386_ VGND VGND VPWR VPWR _1393_ sky130_fd_sc_hd__mux2_1
Xhold110 ram\[5\]\[0\] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dlygate4sd3_1
X_2778_ net162 _1325_ _1349_ VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold132 ram\[17\]\[4\] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 ram\[55\]\[2\] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 ram\[24\]\[5\] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__dlygate4sd3_1
X_1729_ _0533_ addr_reg\[1\] _0531_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__mux2_1
Xhold154 ram\[0\]\[1\] VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 ram\[59\]\[0\] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 ram\[21\]\[4\] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 ram\[52\]\[4\] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 ram\[15\]\[7\] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3750_ clknet_leaf_20_clk _0312_ VGND VGND VPWR VPWR ram\[43\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2701_ _1310_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3681_ clknet_leaf_14_clk _0243_ VGND VGND VPWR VPWR ram\[34\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2632_ net39 _1196_ _1267_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2563_ _1236_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2494_ net43 _1198_ _1184_ VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__mux2_1
X_3115_ net10 VGND VGND VPWR VPWR _1544_ sky130_fd_sc_hd__buf_2
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3046_ _1406_ net180 _1499_ VGND VGND VPWR VPWR _1505_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3948_ clknet_leaf_27_clk _0504_ VGND VGND VPWR VPWR ram\[49\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3879_ clknet_leaf_35_clk _0441_ VGND VGND VPWR VPWR ram\[5\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3802_ clknet_leaf_23_clk _0364_ VGND VGND VPWR VPWR ram\[50\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1994_ _0600_ ram\[60\]\[3\] VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__and2b_1
XFILLER_0_27_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3733_ clknet_leaf_18_clk _0295_ VGND VGND VPWR VPWR ram\[41\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_3664_ clknet_leaf_14_clk _0226_ VGND VGND VPWR VPWR ram\[32\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2615_ _1264_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3595_ clknet_leaf_44_clk _0157_ VGND VGND VPWR VPWR ram\[24\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2546_ _1227_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__clkbuf_1
X_2477_ _1187_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3029_ _1495_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2400_ net70 _1058_ _1139_ VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__mux2_1
X_3380_ _1687_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__clkbuf_1
X_2331_ _1101_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__clkbuf_1
X_2262_ _1050_ _1053_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__nor2_4
XFILLER_0_79_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2193_ ram\[32\]\[6\] ram\[33\]\[6\] ram\[34\]\[6\] ram\[35\]\[6\] _0629_ _0550_
+ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__mux4_1
XFILLER_0_62_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3716_ clknet_leaf_41_clk _0278_ VGND VGND VPWR VPWR ram\[3\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1977_ _0560_ _0773_ _0564_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__o21a_1
X_3647_ clknet_leaf_8_clk _0209_ VGND VGND VPWR VPWR ram\[30\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3578_ clknet_leaf_4_clk _0140_ VGND VGND VPWR VPWR ram\[22\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2529_ _1218_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__clkbuf_1
Xhold14 ram\[15\]\[1\] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold25 ram\[37\]\[6\] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 ram\[34\]\[7\] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 ram\[12\]\[2\] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 ram\[34\]\[6\] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 ram\[44\]\[5\] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2880_ _1414_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__clkbuf_1
X_1900_ ram\[16\]\[1\] ram\[17\]\[1\] ram\[18\]\[1\] ram\[19\]\[1\] _0588_ _0634_
+ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_25_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1831_ _0628_ _0630_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1762_ ram\[42\]\[0\] ram\[43\]\[0\] _0561_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold506 ram\[49\]\[2\] VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__dlygate4sd3_1
X_3501_ clknet_leaf_10_clk _0063_ VGND VGND VPWR VPWR ram\[12\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3432_ net310 net12 _1709_ VGND VGND VPWR VPWR _1715_ sky130_fd_sc_hd__mux2_1
X_3363_ _1678_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__clkbuf_1
X_3294_ _1546_ net439 _1637_ VGND VGND VPWR VPWR _1642_ sky130_fd_sc_hd__mux2_1
X_2314_ _1089_ net5 _0540_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__or3_1
X_2245_ _1035_ _1036_ _1037_ _0934_ _0944_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__o221a_1
X_2176_ ram\[54\]\[6\] ram\[55\]\[6\] _0593_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_69_Left_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_78_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2030_ _0554_ _0825_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_65_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2932_ _1443_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_42_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_57_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2863_ _1403_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__clkbuf_1
X_1814_ _0549_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__clkbuf_4
X_2794_ _1364_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__clkbuf_1
X_1745_ _0544_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__clkbuf_4
Xhold303 ram\[20\]\[6\] VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 ram\[30\]\[6\] VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 ram\[8\]\[6\] VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 ram\[24\]\[3\] VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 ram\[1\]\[7\] VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 ram\[10\]\[0\] VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 ram\[43\]\[3\] VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__dlygate4sd3_1
X_3415_ _1064_ net527 _1700_ VGND VGND VPWR VPWR _1706_ sky130_fd_sc_hd__mux2_1
X_3346_ _1669_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__clkbuf_1
X_3277_ _1546_ net492 _1628_ VGND VGND VPWR VPWR _1633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2228_ _0554_ _1020_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__or2_1
X_2159_ _0546_ _0948_ _0950_ _0952_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_36_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_33_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_70_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3200_ _1094_ _1591_ VGND VGND VPWR VPWR _1592_ sky130_fd_sc_hd__nor2b_4
XFILLER_0_38_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3131_ _1537_ net450 _1554_ VGND VGND VPWR VPWR _1555_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3062_ _1514_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__clkbuf_1
X_2013_ _0806_ _0808_ _0809_ _0564_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_15_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_2
X_3964_ clknet_leaf_16_clk _0520_ VGND VGND VPWR VPWR ram\[39\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2915_ net328 _1315_ _1432_ VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__mux2_1
X_3895_ clknet_leaf_30_clk _0457_ VGND VGND VPWR VPWR ram\[61\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2846_ _1392_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold100 ram\[22\]\[2\] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dlygate4sd3_1
X_2777_ _1355_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__clkbuf_1
Xhold133 ram\[4\]\[5\] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 ram\[24\]\[0\] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dlygate4sd3_1
X_1728_ net2 VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__buf_2
Xhold111 ram\[29\]\[2\] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 ram\[31\]\[2\] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 ram\[43\]\[7\] VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 ram\[10\]\[7\] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 ram\[42\]\[5\] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 ram\[1\]\[1\] VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 ram\[22\]\[3\] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__dlygate4sd3_1
X_3329_ _1660_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2700_ net102 _1196_ _1303_ VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3680_ clknet_leaf_14_clk _0242_ VGND VGND VPWR VPWR ram\[34\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2631_ _1273_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2562_ net326 _1196_ _1229_ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__mux2_1
X_2493_ net14 VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_4_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_2
X_3114_ _1543_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_38_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3045_ _1504_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3947_ clknet_leaf_30_clk _0503_ VGND VGND VPWR VPWR ram\[49\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3878_ clknet_leaf_35_clk _0440_ VGND VGND VPWR VPWR ram\[5\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2829_ _1383_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3801_ clknet_leaf_37_clk _0363_ VGND VGND VPWR VPWR ram\[4\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1993_ _0785_ _0789_ _0598_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__o21ba_1
X_3732_ clknet_leaf_17_clk _0294_ VGND VGND VPWR VPWR ram\[41\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_41_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3663_ clknet_leaf_16_clk _0225_ VGND VGND VPWR VPWR ram\[32\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2614_ net287 _1196_ _1257_ VGND VGND VPWR VPWR _1264_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3594_ clknet_leaf_2_clk _0156_ VGND VGND VPWR VPWR ram\[24\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2545_ net158 _1196_ _1220_ VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__mux2_1
X_2476_ net276 _1186_ _1184_ VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_50_Left_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3028_ _1406_ net139 _1489_ VGND VGND VPWR VPWR _1495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2330_ net51 _1064_ _1095_ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__mux2_1
X_2261_ _1052_ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__clkbuf_8
X_2192_ _0983_ _0984_ _0985_ _0934_ _0585_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__o221a_1
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1976_ ram\[42\]\[3\] ram\[43\]\[3\] _0561_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3715_ clknet_leaf_44_clk _0277_ VGND VGND VPWR VPWR ram\[3\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3646_ clknet_leaf_7_clk _0208_ VGND VGND VPWR VPWR ram\[30\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3577_ clknet_leaf_3_clk _0139_ VGND VGND VPWR VPWR ram\[21\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2528_ net96 _1196_ _1211_ VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold26 ram\[20\]\[2\] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 ram\[48\]\[7\] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 ram\[15\]\[2\] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dlygate4sd3_1
X_2459_ net380 _1060_ _1172_ VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__mux2_1
Xhold48 ram\[54\]\[2\] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 ram\[1\]\[5\] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_7_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1830_ ram\[20\]\[0\] ram\[21\]\[0\] _0629_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1761_ _0555_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__clkbuf_8
X_3500_ clknet_leaf_9_clk _0062_ VGND VGND VPWR VPWR ram\[12\]\[2\] sky130_fd_sc_hd__dfxtp_1
Xhold507 ram\[11\]\[4\] VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__dlygate4sd3_1
X_3431_ _1714_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__clkbuf_1
X_3362_ _1062_ net364 _1673_ VGND VGND VPWR VPWR _1678_ sky130_fd_sc_hd__mux2_1
X_2313_ net4 VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__inv_2
X_3293_ _1641_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__clkbuf_1
X_2244_ ram\[42\]\[7\] ram\[43\]\[7\] _0733_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2175_ _0590_ ram\[53\]\[6\] _0591_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1959_ ram\[12\]\[2\] ram\[13\]\[2\] ram\[14\]\[2\] ram\[15\]\[2\] _0638_ _0624_
+ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__mux4_1
X_3629_ clknet_leaf_7_clk _0191_ VGND VGND VPWR VPWR ram\[28\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput16 net16 VGND VGND VPWR VPWR q[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2931_ _1395_ net47 _1442_ VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_2862_ _1402_ net95 _1396_ VGND VGND VPWR VPWR _1403_ sky130_fd_sc_hd__mux2_1
X_1813_ _0584_ _0599_ _0612_ _0005_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__o31a_1
X_2793_ net55 _1323_ _1358_ VGND VGND VPWR VPWR _1364_ sky130_fd_sc_hd__mux2_1
X_1744_ _0002_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__clkbuf_4
Xhold326 ram\[33\]\[2\] VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold304 ram\[7\]\[6\] VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 ram\[20\]\[1\] VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 ram\[34\]\[3\] VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__dlygate4sd3_1
X_3414_ _1705_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__clkbuf_1
Xhold337 ram\[2\]\[5\] VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold359 ram\[29\]\[7\] VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3345_ net150 net11 _1664_ VGND VGND VPWR VPWR _1669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3276_ _1632_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__clkbuf_1
X_2227_ ram\[56\]\[7\] ram\[57\]\[7\] _0593_ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2158_ _0595_ _0951_ _0944_ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2089_ _0568_ ram\[36\]\[5\] VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_36_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3130_ _1470_ _1509_ VGND VGND VPWR VPWR _1554_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_78_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3061_ net323 _1319_ _1510_ VGND VGND VPWR VPWR _1514_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2012_ ram\[16\]\[3\] ram\[17\]\[3\] ram\[18\]\[3\] ram\[19\]\[3\] _0561_ _0634_
+ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__mux4_2
XFILLER_0_54_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3963_ clknet_leaf_15_clk _0519_ VGND VGND VPWR VPWR ram\[39\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_3894_ clknet_leaf_32_clk _0456_ VGND VGND VPWR VPWR ram\[61\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2914_ _1433_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__clkbuf_1
X_2845_ net201 _1323_ _1386_ VGND VGND VPWR VPWR _1392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold101 ram\[63\]\[2\] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dlygate4sd3_1
X_2776_ net126 _1323_ _1349_ VGND VGND VPWR VPWR _1355_ sky130_fd_sc_hd__mux2_1
Xhold123 ram\[0\]\[2\] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 ram\[3\]\[2\] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dlygate4sd3_1
X_1727_ _0532_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__clkbuf_1
Xhold134 ram\[44\]\[6\] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 ram\[58\]\[3\] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 ram\[23\]\[1\] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 ram\[32\]\[0\] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 ram\[36\]\[5\] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 ram\[14\]\[1\] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__dlygate4sd3_1
X_3328_ net195 net11 _1655_ VGND VGND VPWR VPWR _1660_ sky130_fd_sc_hd__mux2_1
X_3259_ _1623_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_75_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2630_ net166 _1194_ _1267_ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__mux2_1
X_2561_ _1235_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2492_ _1197_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__clkbuf_1
X_3113_ _1542_ net521 _1538_ VGND VGND VPWR VPWR _1543_ sky130_fd_sc_hd__mux2_1
X_3044_ _1404_ net509 _1499_ VGND VGND VPWR VPWR _1504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3946_ clknet_leaf_36_clk _0502_ VGND VGND VPWR VPWR ram\[49\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3877_ clknet_leaf_40_clk _0439_ VGND VGND VPWR VPWR ram\[5\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2828_ _1083_ net245 _1377_ VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__mux2_1
X_2759_ _1085_ net377 _1338_ VGND VGND VPWR VPWR _1345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3800_ clknet_leaf_37_clk _0362_ VGND VGND VPWR VPWR ram\[4\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_43_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3731_ clknet_leaf_17_clk _0293_ VGND VGND VPWR VPWR ram\[41\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_1992_ _0786_ _0787_ _0788_ _0595_ _0596_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__o221a_1
XFILLER_0_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3662_ clknet_leaf_12_clk _0224_ VGND VGND VPWR VPWR ram\[32\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2613_ _1263_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__clkbuf_1
X_3593_ clknet_leaf_4_clk _0155_ VGND VGND VPWR VPWR ram\[23\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2544_ _1226_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2475_ net8 VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__buf_2
XFILLER_0_76_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3027_ _1494_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3929_ clknet_leaf_36_clk _0485_ VGND VGND VPWR VPWR ram\[63\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2260_ _1051_ _0537_ net5 net6 VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2191_ ram\[38\]\[6\] ram\[39\]\[6\] _0733_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1975_ _0554_ _0771_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__or2_1
X_3714_ clknet_leaf_42_clk _0276_ VGND VGND VPWR VPWR ram\[3\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_3645_ clknet_leaf_7_clk _0207_ VGND VGND VPWR VPWR ram\[30\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3576_ clknet_leaf_3_clk _0138_ VGND VGND VPWR VPWR ram\[21\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2527_ _1217_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2458_ _1175_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_3_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold16 ram\[24\]\[6\] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 ram\[48\]\[6\] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 ram\[23\]\[7\] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 ram\[17\]\[6\] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dlygate4sd3_1
X_2389_ _1085_ net435 _1128_ VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1760_ _0559_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__clkbuf_4
Xhold508 ram\[61\]\[0\] VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3430_ net191 net11 _1709_ VGND VGND VPWR VPWR _1714_ sky130_fd_sc_hd__mux2_1
X_3361_ _1677_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2312_ _1088_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__clkbuf_1
X_3292_ _1544_ net459 _1637_ VGND VGND VPWR VPWR _1641_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2243_ _0600_ ram\[41\]\[7\] _0577_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__a21o_1
X_2174_ _0623_ ram\[52\]\[6\] VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1958_ _0752_ _0754_ _0755_ _0564_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__a22o_1
X_1889_ _0584_ _0680_ _0687_ _0005_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__o31a_1
XFILLER_0_3_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3628_ clknet_leaf_6_clk _0190_ VGND VGND VPWR VPWR ram\[28\]\[2\] sky130_fd_sc_hd__dfxtp_1
Xoutput17 net17 VGND VGND VPWR VPWR q[1] sky130_fd_sc_hd__clkbuf_4
X_3559_ clknet_leaf_40_clk _0121_ VGND VGND VPWR VPWR ram\[1\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2930_ _1441_ _1431_ VGND VGND VPWR VPWR _1442_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_73_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2861_ net10 VGND VGND VPWR VPWR _1402_ sky130_fd_sc_hd__clkbuf_4
X_1812_ _0607_ _0610_ _0611_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2792_ _1363_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__clkbuf_1
X_1743_ _0542_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__clkbuf_4
Xhold305 ram\[40\]\[1\] VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 ram\[51\]\[1\] VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__dlygate4sd3_1
X_3413_ _1062_ net281 _1700_ VGND VGND VPWR VPWR _1705_ sky130_fd_sc_hd__mux2_1
Xhold327 ram\[4\]\[3\] VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold338 ram\[53\]\[1\] VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold349 ram\[55\]\[7\] VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3344_ _1668_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__clkbuf_1
X_3275_ _1544_ net300 _1628_ VGND VGND VPWR VPWR _1632_ sky130_fd_sc_hd__mux2_1
X_2226_ ram\[60\]\[7\] ram\[61\]\[7\] ram\[62\]\[7\] ram\[63\]\[7\] _0548_ _0551_
+ VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2157_ ram\[10\]\[6\] ram\[11\]\[6\] _0593_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__mux2_1
X_2088_ _0546_ _0878_ _0880_ _0882_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3060_ _1513_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__clkbuf_1
X_2011_ _0559_ _0807_ _0544_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3962_ clknet_leaf_16_clk _0518_ VGND VGND VPWR VPWR ram\[39\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3893_ clknet_leaf_31_clk _0455_ VGND VGND VPWR VPWR ram\[61\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2913_ net125 _1312_ _1432_ VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__mux2_1
X_2844_ _1391_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__clkbuf_1
X_2775_ _1354_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__clkbuf_1
Xhold135 ram\[1\]\[6\] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 ram\[1\]\[2\] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 ram\[63\]\[5\] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dlygate4sd3_1
X_1726_ _0530_ net463 _0531_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__mux2_1
Xhold102 ram\[40\]\[0\] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 ram\[20\]\[7\] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 ram\[47\]\[5\] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 ram\[39\]\[4\] VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 ram\[33\]\[6\] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__dlygate4sd3_1
X_3327_ _1659_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__clkbuf_1
X_3258_ net298 net10 _1619_ VGND VGND VPWR VPWR _1623_ sky130_fd_sc_hd__mux2_1
X_3189_ _1585_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__clkbuf_1
X_2209_ _0999_ _1000_ _1001_ _0934_ _0944_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_49_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2560_ net311 _1194_ _1229_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__mux2_1
X_2491_ net34 _1196_ _1184_ VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3112_ net9 VGND VGND VPWR VPWR _1542_ sky130_fd_sc_hd__buf_2
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3043_ _1503_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_46_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3945_ clknet_leaf_27_clk _0501_ VGND VGND VPWR VPWR ram\[49\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3876_ clknet_leaf_35_clk _0438_ VGND VGND VPWR VPWR ram\[5\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2827_ _1382_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__clkbuf_1
X_2758_ _1344_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2689_ _1304_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_1_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1991_ ram\[50\]\[3\] ram\[51\]\[3\] _0733_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3730_ clknet_leaf_18_clk _0292_ VGND VGND VPWR VPWR ram\[41\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3661_ clknet_leaf_16_clk _0223_ VGND VGND VPWR VPWR ram\[32\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_3592_ clknet_leaf_2_clk _0154_ VGND VGND VPWR VPWR ram\[23\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2612_ net346 _1194_ _1257_ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2543_ net82 _1194_ _1220_ VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2474_ _1185_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3026_ _1404_ net485 _1489_ VGND VGND VPWR VPWR _1494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3928_ clknet_leaf_33_clk _0484_ VGND VGND VPWR VPWR ram\[63\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3859_ clknet_leaf_36_clk _0421_ VGND VGND VPWR VPWR ram\[57\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2190_ _0568_ ram\[37\]\[6\] _0577_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1974_ ram\[40\]\[3\] ram\[41\]\[3\] _0556_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__mux2_1
X_3713_ clknet_leaf_15_clk _0275_ VGND VGND VPWR VPWR ram\[38\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3644_ clknet_leaf_7_clk _0206_ VGND VGND VPWR VPWR ram\[30\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3575_ clknet_leaf_1_clk _0137_ VGND VGND VPWR VPWR ram\[21\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2526_ net425 _1194_ _1211_ VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2457_ net60 _1058_ _1172_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold28 ram\[8\]\[5\] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 ram\[13\]\[2\] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold39 ram\[23\]\[0\] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dlygate4sd3_1
X_2388_ _1134_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_54_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3009_ _1404_ net428 _1480_ VGND VGND VPWR VPWR _1485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3360_ _1060_ net458 _1673_ VGND VGND VPWR VPWR _1677_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_29_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2311_ _1087_ net382 _1073_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__mux2_1
X_3291_ _1640_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2242_ _0651_ ram\[40\]\[7\] VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__and2b_1
X_2173_ _0546_ _0962_ _0964_ _0966_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1957_ ram\[16\]\[2\] ram\[17\]\[2\] ram\[18\]\[2\] ram\[19\]\[2\] _0561_ _0634_
+ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__mux4_2
XFILLER_0_7_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1888_ _0684_ _0686_ _0611_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3627_ clknet_leaf_0_clk _0189_ VGND VGND VPWR VPWR ram\[28\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_3558_ clknet_leaf_41_clk _0120_ VGND VGND VPWR VPWR ram\[1\]\[4\] sky130_fd_sc_hd__dfxtp_1
Xoutput18 net18 VGND VGND VPWR VPWR q[2] sky130_fd_sc_hd__clkbuf_4
X_2509_ net525 _1194_ _1202_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__mux2_1
X_3489_ clknet_leaf_13_clk _0051_ VGND VGND VPWR VPWR ram\[10\]\[7\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_36_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_27_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_69_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2860_ _1401_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_73_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1811_ _0003_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__buf_4
XFILLER_0_72_327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2791_ net330 _1321_ _1358_ VGND VGND VPWR VPWR _1363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1742_ _0003_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__clkbuf_4
Xhold317 ram\[41\]\[1\] VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold306 ram\[22\]\[6\] VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__dlygate4sd3_1
X_3412_ _1704_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__clkbuf_1
Xhold339 ram\[49\]\[5\] VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 ram\[21\]\[5\] VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3343_ net171 net10 _1664_ VGND VGND VPWR VPWR _1668_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3274_ _1631_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__clkbuf_1
X_2225_ _0611_ _1010_ _1017_ _0581_ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__a211o_1
X_2156_ _0554_ _0949_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_64_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2087_ _0560_ _0881_ _0564_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_18_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_75_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2989_ _1474_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2010_ ram\[22\]\[3\] ram\[23\]\[3\] _0608_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__mux2_1
X_3961_ clknet_leaf_16_clk _0517_ VGND VGND VPWR VPWR ram\[39\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2912_ _1094_ _1431_ VGND VGND VPWR VPWR _1432_ sky130_fd_sc_hd__nor2b_4
X_3892_ clknet_leaf_32_clk _0454_ VGND VGND VPWR VPWR ram\[61\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2843_ net93 _1321_ _1386_ VGND VGND VPWR VPWR _1391_ sky130_fd_sc_hd__mux2_1
X_2774_ net97 _1321_ _1349_ VGND VGND VPWR VPWR _1354_ sky130_fd_sc_hd__mux2_1
X_1725_ net15 VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold114 ram\[0\]\[0\] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 ram\[1\]\[4\] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 ram\[32\]\[5\] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 ram\[6\]\[5\] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 ram\[19\]\[3\] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_2
Xhold147 ram\[8\]\[0\] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 ram\[3\]\[5\] VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3326_ net107 net10 _1655_ VGND VGND VPWR VPWR _1659_ sky130_fd_sc_hd__mux2_1
X_3257_ _1622_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__clkbuf_1
X_2208_ ram\[18\]\[7\] ram\[19\]\[7\] _0654_ VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__mux2_1
X_3188_ _1544_ net442 _1581_ VGND VGND VPWR VPWR _1585_ sky130_fd_sc_hd__mux2_1
X_2139_ _0551_ _0932_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_49_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2490_ net13 VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__buf_2
XFILLER_0_50_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3111_ _1541_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__clkbuf_1
X_3042_ _1402_ net526 _1499_ VGND VGND VPWR VPWR _1503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3944_ clknet_leaf_27_clk _0500_ VGND VGND VPWR VPWR ram\[49\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3875_ clknet_leaf_39_clk _0437_ VGND VGND VPWR VPWR ram\[5\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2826_ _1081_ net502 _1377_ VGND VGND VPWR VPWR _1382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2757_ _1083_ net443 _1338_ VGND VGND VPWR VPWR _1344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2688_ net118 _1181_ _1303_ VGND VGND VPWR VPWR _1304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3309_ _1544_ net233 _1646_ VGND VGND VPWR VPWR _1650_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1990_ _0590_ ram\[49\]\[3\] _0591_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_43_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3660_ clknet_leaf_11_clk _0222_ VGND VGND VPWR VPWR ram\[32\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3591_ clknet_leaf_1_clk _0153_ VGND VGND VPWR VPWR ram\[23\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2611_ _1262_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__clkbuf_1
X_2542_ _1225_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__clkbuf_1
X_2473_ net203 _1181_ _1184_ VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3025_ _1493_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__clkbuf_1
X_3927_ clknet_leaf_37_clk _0483_ VGND VGND VPWR VPWR ram\[6\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3858_ clknet_leaf_36_clk _0420_ VGND VGND VPWR VPWR ram\[57\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_3789_ clknet_leaf_36_clk _0351_ VGND VGND VPWR VPWR ram\[48\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2809_ _1372_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1973_ ram\[44\]\[3\] ram\[45\]\[3\] ram\[46\]\[3\] ram\[47\]\[3\] _0548_ _0551_
+ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3712_ clknet_leaf_25_clk _0274_ VGND VGND VPWR VPWR ram\[38\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3643_ clknet_leaf_0_clk _0205_ VGND VGND VPWR VPWR ram\[30\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3574_ clknet_leaf_6_clk _0136_ VGND VGND VPWR VPWR ram\[21\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2525_ _1216_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__clkbuf_1
X_2456_ _1174_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__clkbuf_1
Xhold18 ram\[18\]\[7\] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 ram\[8\]\[3\] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2387_ _1083_ net303 _1128_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3008_ _1484_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3290_ _1542_ net424 _1637_ VGND VGND VPWR VPWR _1640_ sky130_fd_sc_hd__mux2_1
X_2310_ net14 VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__buf_2
X_2241_ _0545_ _1033_ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2172_ _0560_ _0965_ _0575_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_51_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1956_ _0559_ _0753_ _0544_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1887_ _0575_ _0685_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3626_ clknet_leaf_5_clk _0188_ VGND VGND VPWR VPWR ram\[28\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_3557_ clknet_leaf_40_clk _0119_ VGND VGND VPWR VPWR ram\[1\]\[3\] sky130_fd_sc_hd__dfxtp_1
Xoutput19 net19 VGND VGND VPWR VPWR q[3] sky130_fd_sc_hd__clkbuf_4
X_2508_ _1207_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__clkbuf_1
X_3488_ clknet_leaf_13_clk _0050_ VGND VGND VPWR VPWR ram\[10\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2439_ _1077_ net109 _1162_ VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1810_ _0575_ _0609_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__and2_1
X_2790_ _1362_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1741_ _0541_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold307 ram\[33\]\[4\] VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__dlygate4sd3_1
X_3411_ _1060_ net181 _1700_ VGND VGND VPWR VPWR _1704_ sky130_fd_sc_hd__mux2_1
Xhold318 ram\[6\]\[6\] VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 ram\[34\]\[4\] VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__dlygate4sd3_1
X_3342_ _1667_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3273_ _1542_ net103 _1628_ VGND VGND VPWR VPWR _1631_ sky130_fd_sc_hd__mux2_1
X_2224_ _1014_ _1016_ _0003_ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__o21ba_1
X_2155_ ram\[8\]\[6\] ram\[9\]\[6\] _0733_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__mux2_1
X_2086_ ram\[42\]\[5\] ram\[43\]\[5\] _0651_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2988_ _1400_ net523 _1471_ VGND VGND VPWR VPWR _1474_ sky130_fd_sc_hd__mux2_1
X_1939_ _0600_ ram\[60\]\[2\] VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__and2b_1
X_3609_ clknet_leaf_38_clk _0171_ VGND VGND VPWR VPWR ram\[25\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Left_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Left_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3960_ clknet_leaf_16_clk _0516_ VGND VGND VPWR VPWR ram\[39\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2911_ _1430_ VGND VGND VPWR VPWR _1431_ sky130_fd_sc_hd__buf_6
X_3891_ clknet_leaf_30_clk _0453_ VGND VGND VPWR VPWR ram\[61\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_75_Left_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2842_ _1390_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2773_ _1353_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1724_ net1 VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold115 ram\[17\]\[2\] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 ram\[26\]\[3\] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 ram\[22\]\[7\] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 ram\[7\]\[1\] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold148 ram\[6\]\[3\] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 ram\[5\]\[5\] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3325_ _1658_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__clkbuf_1
X_3256_ net227 net9 _1619_ VGND VGND VPWR VPWR _1622_ sky130_fd_sc_hd__mux2_1
X_2207_ _0588_ ram\[17\]\[7\] _0553_ VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__a21o_1
X_3187_ _1584_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2138_ ram\[28\]\[6\] ram\[29\]\[6\] _0654_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2069_ ram\[12\]\[4\] ram\[13\]\[4\] ram\[14\]\[4\] ram\[15\]\[4\] _0600_ _0624_
+ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__mux4_1
XFILLER_0_8_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3110_ _1540_ net339 _1538_ VGND VGND VPWR VPWR _1541_ sky130_fd_sc_hd__mux2_1
X_3041_ _1502_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__clkbuf_1
X_3943_ clknet_leaf_27_clk _0499_ VGND VGND VPWR VPWR ram\[59\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3874_ clknet_leaf_40_clk _0436_ VGND VGND VPWR VPWR ram\[5\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2825_ _1381_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2756_ _1343_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__clkbuf_1
X_2687_ _1266_ _1137_ VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__nor2_4
XFILLER_0_41_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3308_ _1649_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__clkbuf_1
X_3239_ _1542_ net250 _1610_ VGND VGND VPWR VPWR _1613_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold490 ram\[24\]\[2\] VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3590_ clknet_leaf_5_clk _0152_ VGND VGND VPWR VPWR ram\[23\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2610_ net113 _1192_ _1257_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__mux2_1
X_2541_ net148 _1192_ _1220_ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2472_ _1094_ _1183_ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__nor2_4
XFILLER_0_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3024_ _1402_ net514 _1489_ VGND VGND VPWR VPWR _1493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3926_ clknet_leaf_37_clk _0482_ VGND VGND VPWR VPWR ram\[6\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3857_ clknet_leaf_27_clk _0419_ VGND VGND VPWR VPWR ram\[56\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3788_ clknet_leaf_36_clk _0350_ VGND VGND VPWR VPWR ram\[48\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2808_ net352 _1321_ _1367_ VGND VGND VPWR VPWR _1372_ sky130_fd_sc_hd__mux2_1
X_2739_ _1334_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1972_ _0727_ _0744_ _0769_ _0659_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__a22o_1
X_3711_ clknet_leaf_15_clk _0273_ VGND VGND VPWR VPWR ram\[38\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3642_ clknet_leaf_7_clk _0204_ VGND VGND VPWR VPWR ram\[30\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3573_ clknet_leaf_6_clk _0135_ VGND VGND VPWR VPWR ram\[21\]\[3\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2524_ net373 _1192_ _1211_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__mux2_1
X_2455_ net37 _1056_ _1172_ VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__mux2_1
Xhold19 ram\[12\]\[1\] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlygate4sd3_1
X_2386_ _1133_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_3_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3007_ _1402_ net481 _1480_ VGND VGND VPWR VPWR _1484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3909_ clknet_leaf_14_clk _0009_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_34_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2240_ ram\[44\]\[7\] ram\[45\]\[7\] ram\[46\]\[7\] ram\[47\]\[7\] _0567_ _0728_
+ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__mux4_1
X_2171_ ram\[58\]\[6\] ram\[59\]\[6\] _0556_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1955_ ram\[22\]\[2\] ram\[23\]\[2\] _0608_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__mux2_1
X_1886_ ram\[56\]\[1\] ram\[57\]\[1\] ram\[58\]\[1\] ram\[59\]\[1\] _0608_ _0553_
+ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__mux4_1
XFILLER_0_3_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3625_ clknet_leaf_2_clk _0187_ VGND VGND VPWR VPWR ram\[27\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3556_ clknet_leaf_41_clk _0118_ VGND VGND VPWR VPWR ram\[1\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2507_ net155 _1192_ _1202_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__mux2_1
X_3487_ clknet_leaf_5_clk _0049_ VGND VGND VPWR VPWR ram\[10\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2438_ _1164_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__clkbuf_1
X_2369_ _1122_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1740_ _0540_ net24 _0531_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__mux2_1
Xhold308 ram\[7\]\[4\] VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3410_ _1703_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold319 ram\[59\]\[7\] VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__dlygate4sd3_1
X_3341_ net204 net9 _1664_ VGND VGND VPWR VPWR _1667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3272_ _1630_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__clkbuf_1
X_2223_ _0645_ _1015_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__and2_1
X_2154_ ram\[12\]\[6\] ram\[13\]\[6\] ram\[14\]\[6\] ram\[15\]\[6\] _0590_ _0614_
+ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__mux4_1
X_2085_ _0554_ _0879_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_64_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2987_ _1473_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1938_ _0730_ _0735_ _0598_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__o21ba_1
X_1869_ ram\[38\]\[1\] ram\[39\]\[1\] _0556_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__mux2_1
X_3608_ clknet_leaf_2_clk _0170_ VGND VGND VPWR VPWR ram\[25\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3539_ clknet_leaf_44_clk _0101_ VGND VGND VPWR VPWR ram\[17\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2910_ net5 net6 _0537_ VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__and3b_1
X_3890_ clknet_leaf_30_clk _0452_ VGND VGND VPWR VPWR ram\[61\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2841_ net452 _1319_ _1386_ VGND VGND VPWR VPWR _1390_ sky130_fd_sc_hd__mux2_1
X_2772_ net295 _1319_ _1349_ VGND VGND VPWR VPWR _1353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold105 ram\[28\]\[7\] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 ram\[46\]\[5\] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 ram\[6\]\[4\] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 ram\[14\]\[6\] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 ram\[31\]\[4\] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3324_ net231 net9 _1655_ VGND VGND VPWR VPWR _1658_ sky130_fd_sc_hd__mux2_1
X_3255_ _1621_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__clkbuf_1
X_2206_ _0641_ ram\[16\]\[7\] VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__and2b_1
X_3186_ _1542_ net144 _1581_ VGND VGND VPWR VPWR _1584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2137_ _0891_ _0906_ _0931_ _0659_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_49_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2068_ _0860_ _0862_ _0863_ _0564_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3040_ _1400_ net510 _1499_ VGND VGND VPWR VPWR _1502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3942_ clknet_leaf_26_clk _0498_ VGND VGND VPWR VPWR ram\[59\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3873_ clknet_leaf_27_clk _0435_ VGND VGND VPWR VPWR ram\[58\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2824_ _1079_ net506 _1377_ VGND VGND VPWR VPWR _1381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2755_ _1081_ net172 _1338_ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__mux2_1
X_2686_ _1302_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3307_ _1542_ net418 _1646_ VGND VGND VPWR VPWR _1649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3238_ _1612_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__clkbuf_1
X_3169_ _1542_ net71 _1572_ VGND VGND VPWR VPWR _1575_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold480 ram\[52\]\[2\] VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold491 ram\[46\]\[3\] VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_43_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2540_ _1224_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__clkbuf_1
X_2471_ _1182_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__buf_4
X_3023_ _1492_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3925_ clknet_leaf_39_clk _0481_ VGND VGND VPWR VPWR ram\[6\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_446 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3856_ clknet_leaf_27_clk _0418_ VGND VGND VPWR VPWR ram\[56\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2807_ _1371_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__clkbuf_1
X_3787_ clknet_leaf_27_clk _0349_ VGND VGND VPWR VPWR ram\[48\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2738_ _1081_ net265 _1329_ VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__mux2_1
X_2669_ _1293_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1971_ _0750_ _0756_ _0762_ _0768_ _0004_ _0611_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__mux4_1
X_3710_ clknet_leaf_15_clk _0272_ VGND VGND VPWR VPWR ram\[38\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3641_ clknet_leaf_37_clk _0203_ VGND VGND VPWR VPWR ram\[2\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3572_ clknet_leaf_6_clk _0134_ VGND VGND VPWR VPWR ram\[21\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2523_ _1215_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2454_ _1173_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__clkbuf_1
X_2385_ _1081_ net530 _1128_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__mux2_1
Xinput1 addr[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XFILLER_0_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3006_ _1483_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3908_ clknet_leaf_26_clk _0008_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3839_ clknet_leaf_30_clk _0401_ VGND VGND VPWR VPWR ram\[54\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_17_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2170_ _0554_ _0963_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1954_ _0628_ _0751_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__or2_1
X_1885_ _0681_ _0682_ _0683_ _0606_ _0573_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__o221a_1
X_3624_ clknet_leaf_2_clk _0186_ VGND VGND VPWR VPWR ram\[27\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3555_ clknet_leaf_2_clk _0117_ VGND VGND VPWR VPWR ram\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2506_ _1206_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__clkbuf_1
X_3486_ clknet_leaf_10_clk _0048_ VGND VGND VPWR VPWR ram\[10\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2437_ _1075_ net212 _1162_ VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2368_ net242 _1066_ _1115_ VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__mux2_1
X_2299_ _1079_ net219 _1073_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold309 ram\[39\]\[7\] VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3340_ _1666_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3271_ _1540_ net478 _1628_ VGND VGND VPWR VPWR _1630_ sky130_fd_sc_hd__mux2_1
X_2222_ ram\[0\]\[7\] ram\[1\]\[7\] ram\[2\]\[7\] ram\[3\]\[7\] _0547_ _0728_ VGND
+ VGND VPWR VPWR _1015_ sky130_fd_sc_hd__mux4_1
X_2153_ _0611_ _0938_ _0946_ _0584_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2084_ ram\[40\]\[5\] ram\[41\]\[5\] _0556_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2986_ _1398_ net471 _1471_ VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__mux2_1
X_1937_ _0731_ _0732_ _0734_ _0595_ _0596_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1868_ _0548_ ram\[37\]\[1\] _0570_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__a21o_1
X_3607_ clknet_leaf_44_clk _0169_ VGND VGND VPWR VPWR ram\[25\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_3538_ clknet_leaf_43_clk _0100_ VGND VGND VPWR VPWR ram\[17\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_1799_ _0587_ _0597_ _0598_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_12_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3469_ clknet_leaf_12_clk _0031_ VGND VGND VPWR VPWR ram\[8\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2840_ _1389_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__clkbuf_1
X_2771_ _1352_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold117 ram\[26\]\[1\] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold106 ram\[15\]\[4\] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 ram\[4\]\[2\] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold139 ram\[32\]\[6\] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__dlygate4sd3_1
X_3323_ _1657_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__clkbuf_1
X_3254_ net154 net8 _1619_ VGND VGND VPWR VPWR _1621_ sky130_fd_sc_hd__mux2_1
X_2205_ _0621_ _0997_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__and2_1
X_3185_ _1583_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__clkbuf_1
X_2136_ _0912_ _0918_ _0924_ _0930_ _0611_ _0584_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__mux4_1
X_2067_ ram\[16\]\[4\] ram\[17\]\[4\] ram\[18\]\[4\] ram\[19\]\[4\] _0561_ _0634_
+ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_49_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2969_ _1463_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3941_ clknet_leaf_36_clk _0497_ VGND VGND VPWR VPWR ram\[59\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3872_ clknet_leaf_26_clk _0434_ VGND VGND VPWR VPWR ram\[58\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2823_ _1380_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__clkbuf_1
X_2754_ _1342_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2685_ _1087_ net391 _1294_ VGND VGND VPWR VPWR _1302_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3306_ _1648_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__clkbuf_1
X_3237_ _1540_ net480 _1610_ VGND VGND VPWR VPWR _1612_ sky130_fd_sc_hd__mux2_1
X_3168_ _1574_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__clkbuf_1
X_2119_ _0628_ _0913_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__or2_1
X_3099_ _1406_ ram\[50\]\[5\] _1528_ VGND VGND VPWR VPWR _1534_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold470 ram\[50\]\[6\] VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 ram\[9\]\[1\] VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 ram\[61\]\[5\] VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_43_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2470_ _0537_ _1124_ _0540_ VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__or3_1
X_3022_ _1400_ net444 _1489_ VGND VGND VPWR VPWR _1492_ sky130_fd_sc_hd__mux2_1
X_3924_ clknet_leaf_41_clk _0480_ VGND VGND VPWR VPWR ram\[6\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3855_ clknet_leaf_33_clk _0417_ VGND VGND VPWR VPWR ram\[56\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_3786_ clknet_leaf_36_clk _0348_ VGND VGND VPWR VPWR ram\[48\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2806_ net371 _1319_ _1367_ VGND VGND VPWR VPWR _1371_ sky130_fd_sc_hd__mux2_1
X_2737_ _1333_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2668_ net226 _1198_ _1285_ VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2599_ _1087_ net127 _1248_ VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1970_ _0637_ _0763_ _0767_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3640_ clknet_leaf_35_clk _0202_ VGND VGND VPWR VPWR ram\[2\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3571_ clknet_leaf_1_clk _0133_ VGND VGND VPWR VPWR ram\[21\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2522_ net489 _1190_ _1211_ VGND VGND VPWR VPWR _1215_ sky130_fd_sc_hd__mux2_1
X_2453_ net238 _1048_ _1172_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__mux2_1
X_2384_ _1132_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__clkbuf_1
Xinput2 addr[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
X_3005_ _1400_ net501 _1480_ VGND VGND VPWR VPWR _1483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3907_ clknet_leaf_26_clk _0007_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3838_ clknet_leaf_31_clk _0400_ VGND VGND VPWR VPWR ram\[54\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3769_ clknet_leaf_22_clk _0331_ VGND VGND VPWR VPWR ram\[45\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1953_ ram\[20\]\[2\] ram\[21\]\[2\] _0629_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1884_ ram\[62\]\[1\] ram\[63\]\[1\] _0604_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__mux2_1
X_3623_ clknet_leaf_1_clk _0185_ VGND VGND VPWR VPWR ram\[27\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_3554_ clknet_leaf_42_clk _0116_ VGND VGND VPWR VPWR ram\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2505_ net394 _1190_ _1202_ VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__mux2_1
X_3485_ clknet_leaf_11_clk _0047_ VGND VGND VPWR VPWR ram\[10\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2436_ _1163_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2367_ _1121_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__clkbuf_1
X_2298_ net10 VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_67_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3270_ _1629_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2221_ _1011_ _1012_ _1013_ _0934_ _0545_ VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__o221a_1
X_2152_ _0940_ _0945_ _0003_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__o21ba_1
X_2083_ ram\[44\]\[5\] ram\[45\]\[5\] ram\[46\]\[5\] ram\[47\]\[5\] _0548_ _0551_
+ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_64_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2985_ _1472_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__clkbuf_1
X_1936_ ram\[50\]\[2\] ram\[51\]\[2\] _0733_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1867_ _0568_ ram\[36\]\[1\] VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__and2b_1
X_3606_ clknet_leaf_1_clk _0168_ VGND VGND VPWR VPWR ram\[25\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_1798_ _0003_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3537_ clknet_leaf_38_clk _0099_ VGND VGND VPWR VPWR ram\[16\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3468_ clknet_leaf_10_clk _0030_ VGND VGND VPWR VPWR ram\[8\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3399_ _1697_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__clkbuf_1
X_2419_ _1077_ net40 _1150_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2770_ net495 _1317_ _1349_ VGND VGND VPWR VPWR _1352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold107 ram\[20\]\[3\] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 ram\[17\]\[0\] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 ram\[40\]\[7\] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3322_ net504 net8 _1655_ VGND VGND VPWR VPWR _1657_ sky130_fd_sc_hd__mux2_1
X_3253_ _1620_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__clkbuf_1
X_3184_ _1540_ net302 _1581_ VGND VGND VPWR VPWR _1583_ sky130_fd_sc_hd__mux2_1
X_2204_ ram\[20\]\[7\] ram\[21\]\[7\] ram\[22\]\[7\] ram\[23\]\[7\] _0567_ _0728_
+ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_53_Left_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2135_ _0637_ _0925_ _0929_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__a21o_1
X_2066_ _0559_ _0861_ _0544_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_49_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2968_ _1398_ net440 _1461_ VGND VGND VPWR VPWR _1463_ sky130_fd_sc_hd__mux2_1
X_1919_ ram\[42\]\[2\] ram\[43\]\[2\] _0561_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_62_Left_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2899_ _1424_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_71_Left_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_80_Left_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3940_ clknet_leaf_34_clk _0496_ VGND VGND VPWR VPWR ram\[59\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_46_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3871_ clknet_leaf_33_clk _0433_ VGND VGND VPWR VPWR ram\[58\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2822_ _1077_ ram\[35\]\[2\] _1377_ VGND VGND VPWR VPWR _1380_ sky130_fd_sc_hd__mux2_1
X_2753_ _1079_ net345 _1338_ VGND VGND VPWR VPWR _1342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2684_ _1301_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3305_ _1540_ net53 _1646_ VGND VGND VPWR VPWR _1648_ sky130_fd_sc_hd__mux2_1
X_3236_ _1611_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__clkbuf_1
X_3167_ _1540_ net269 _1572_ VGND VGND VPWR VPWR _1574_ sky130_fd_sc_hd__mux2_1
X_2118_ ram\[28\]\[5\] ram\[29\]\[5\] _0629_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__mux2_1
X_3098_ _1533_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__clkbuf_1
X_2049_ _0600_ ram\[60\]\[4\] VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_80_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold471 ram\[63\]\[1\] VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold460 ram\[49\]\[6\] VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 ram\[46\]\[0\] VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 ram\[47\]\[0\] VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3021_ _1491_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3923_ clknet_leaf_40_clk _0479_ VGND VGND VPWR VPWR ram\[6\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3854_ clknet_leaf_34_clk _0416_ VGND VGND VPWR VPWR ram\[56\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2805_ _1370_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3785_ clknet_leaf_22_clk _0347_ VGND VGND VPWR VPWR ram\[47\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2736_ _1079_ net285 _1329_ VGND VGND VPWR VPWR _1333_ sky130_fd_sc_hd__mux2_1
X_2667_ _1292_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2598_ _1255_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3219_ _1602_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold290 ram\[10\]\[3\] VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3570_ clknet_leaf_6_clk _0132_ VGND VGND VPWR VPWR ram\[21\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2521_ _1214_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2452_ _1091_ _1171_ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__nor2_4
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2383_ _1079_ net490 _1128_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__mux2_1
Xinput3 addr[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3004_ _1482_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_19_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3906_ clknet_leaf_37_clk _0006_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_52_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3837_ clknet_leaf_30_clk _0399_ VGND VGND VPWR VPWR ram\[54\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_3768_ clknet_leaf_22_clk _0330_ VGND VGND VPWR VPWR ram\[45\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2719_ _1322_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3699_ clknet_leaf_19_clk _0261_ VGND VGND VPWR VPWR ram\[37\]\[1\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1952_ _0746_ _0748_ _0749_ _0626_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__a22o_1
X_1883_ _0602_ ram\[61\]\[1\] _0570_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__a21o_1
X_3622_ clknet_leaf_0_clk _0184_ VGND VGND VPWR VPWR ram\[27\]\[4\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3553_ clknet_leaf_38_clk _0115_ VGND VGND VPWR VPWR ram\[18\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2504_ _1205_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__clkbuf_1
X_3484_ clknet_leaf_10_clk _0046_ VGND VGND VPWR VPWR ram\[10\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2435_ _1070_ net419 _1162_ VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__mux2_1
X_2366_ net94 _1064_ _1115_ VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2297_ _1078_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2220_ ram\[6\]\[7\] ram\[7\]\[7\] _0654_ VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__mux2_1
X_2151_ _0941_ _0942_ _0943_ _0934_ _0944_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__o221a_1
X_2082_ _0837_ _0852_ _0877_ _0659_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__a22o_1
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2984_ _1395_ net475 _1471_ VGND VGND VPWR VPWR _1472_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1935_ _0555_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__buf_4
XFILLER_0_56_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1866_ _0546_ _0660_ _0662_ _0664_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3605_ clknet_leaf_44_clk _0167_ VGND VGND VPWR VPWR ram\[25\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_1797_ _0589_ _0592_ _0594_ _0595_ _0596_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__o221a_1
X_3536_ clknet_leaf_38_clk _0098_ VGND VGND VPWR VPWR ram\[16\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3467_ clknet_leaf_10_clk _0029_ VGND VGND VPWR VPWR ram\[8\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_3398_ _1064_ net362 _1691_ VGND VGND VPWR VPWR _1697_ sky130_fd_sc_hd__mux2_1
X_2418_ _1152_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__clkbuf_1
X_2349_ net488 _1066_ _1104_ VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold108 ram\[58\]\[4\] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold119 ram\[38\]\[2\] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3321_ _1656_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3252_ net133 net7 _1619_ VGND VGND VPWR VPWR _1620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3183_ _1582_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__clkbuf_1
X_2203_ _0992_ _0994_ _0995_ _0626_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__a22o_1
X_2134_ _0926_ _0927_ _0928_ _0644_ _0645_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__o221a_1
X_2065_ ram\[22\]\[4\] ram\[23\]\[4\] _0608_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2967_ _1462_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__clkbuf_1
X_2898_ net135 _1317_ _1421_ VGND VGND VPWR VPWR _1424_ sky130_fd_sc_hd__mux2_1
X_1918_ _0554_ _0715_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__or2_1
X_1849_ _0555_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__buf_4
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3519_ clknet_leaf_8_clk _0081_ VGND VGND VPWR VPWR ram\[14\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_20_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_50_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3870_ clknet_leaf_34_clk _0432_ VGND VGND VPWR VPWR ram\[58\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2821_ _1379_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2752_ _1341_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_11_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_30_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2683_ _1085_ net449 _1294_ VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__mux2_1
X_3304_ _1647_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__clkbuf_1
X_3235_ _1537_ net423 _1610_ VGND VGND VPWR VPWR _1611_ sky130_fd_sc_hd__mux2_1
X_3166_ _1573_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2117_ _0637_ _0907_ _0911_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__a21o_1
X_3097_ _1404_ ram\[50\]\[4\] _1528_ VGND VGND VPWR VPWR _1533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2048_ _0839_ _0843_ _0598_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_49_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold472 ram\[32\]\[2\] VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 ram\[29\]\[0\] VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold450 ram\[11\]\[1\] VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 ram\[37\]\[1\] VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 ram\[35\]\[3\] VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_0_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_0_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_2
X_3020_ _1398_ net383 _1489_ VGND VGND VPWR VPWR _1491_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3922_ clknet_leaf_41_clk _0478_ VGND VGND VPWR VPWR ram\[6\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3853_ clknet_leaf_34_clk _0415_ VGND VGND VPWR VPWR ram\[56\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2804_ net284 _1317_ _1367_ VGND VGND VPWR VPWR _1370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3784_ clknet_leaf_22_clk _0346_ VGND VGND VPWR VPWR ram\[47\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2735_ _1332_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__clkbuf_1
X_2666_ net260 _1196_ _1285_ VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__mux2_1
X_2597_ _1085_ net329 _1248_ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3218_ _1537_ net479 _1601_ VGND VGND VPWR VPWR _1602_ sky130_fd_sc_hd__mux2_1
X_3149_ _1564_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold280 ram\[11\]\[5\] VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 ram\[60\]\[5\] VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2520_ net336 _1188_ _1211_ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__mux2_1
X_2451_ net15 _1049_ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__nand2_4
X_2382_ _1131_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__clkbuf_1
Xinput4 addr[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dlymetal6s2s_1
X_3003_ _1398_ net470 _1480_ VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3905_ clknet_leaf_28_clk _0467_ VGND VGND VPWR VPWR ram\[62\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3836_ clknet_leaf_31_clk _0398_ VGND VGND VPWR VPWR ram\[54\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3767_ clknet_leaf_21_clk _0329_ VGND VGND VPWR VPWR ram\[45\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2718_ net353 _1321_ _1313_ VGND VGND VPWR VPWR _1322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3698_ clknet_leaf_19_clk _0260_ VGND VGND VPWR VPWR ram\[37\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2649_ net215 _1196_ _1276_ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1951_ ram\[0\]\[2\] ram\[1\]\[2\] ram\[2\]\[2\] ram\[3\]\[2\] _0623_ _0634_ VGND
+ VGND VPWR VPWR _0749_ sky130_fd_sc_hd__mux4_1
X_1882_ _0600_ ram\[60\]\[1\] VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__and2b_1
X_3621_ clknet_leaf_0_clk _0183_ VGND VGND VPWR VPWR ram\[27\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3552_ clknet_leaf_39_clk _0114_ VGND VGND VPWR VPWR ram\[18\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2503_ net138 _1188_ _1202_ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__mux2_1
X_3483_ clknet_leaf_10_clk _0045_ VGND VGND VPWR VPWR ram\[10\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2434_ _1125_ _1161_ VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__nand2_4
X_2365_ _1120_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2296_ _1077_ net134 _1073_ VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3819_ clknet_leaf_29_clk _0381_ VGND VGND VPWR VPWR ram\[52\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2150_ _0563_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__clkbuf_4
X_2081_ _0858_ _0864_ _0870_ _0876_ _0004_ _0611_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2983_ _1470_ _1431_ VGND VGND VPWR VPWR _1471_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_72_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1934_ _0590_ ram\[49\]\[2\] _0591_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1865_ _0560_ _0663_ _0564_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__o21a_1
X_3604_ clknet_leaf_44_clk _0166_ VGND VGND VPWR VPWR ram\[25\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_1796_ _0563_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__buf_2
X_3535_ clknet_leaf_44_clk _0097_ VGND VGND VPWR VPWR ram\[16\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3466_ clknet_leaf_5_clk _0028_ VGND VGND VPWR VPWR ram\[8\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2417_ _1075_ net54 _1150_ VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__mux2_1
X_3397_ _1696_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2348_ _1110_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__clkbuf_1
X_2279_ _1065_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_27_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold109 ram\[36\]\[6\] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3320_ net111 net7 _1655_ VGND VGND VPWR VPWR _1656_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3251_ _1053_ _1072_ VGND VGND VPWR VPWR _1619_ sky130_fd_sc_hd__nor2b_4
X_3182_ _1537_ net405 _1581_ VGND VGND VPWR VPWR _1582_ sky130_fd_sc_hd__mux2_1
X_2202_ ram\[24\]\[7\] ram\[25\]\[7\] ram\[26\]\[7\] ram\[27\]\[7\] _0602_ _0614_
+ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__mux4_1
X_2133_ ram\[10\]\[5\] ram\[11\]\[5\] _0619_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__mux2_1
X_2064_ _0628_ _0859_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2966_ _1395_ net520 _1461_ VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__mux2_1
X_1917_ ram\[40\]\[2\] ram\[41\]\[2\] _0556_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__mux2_1
X_2897_ _1423_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1848_ ram\[28\]\[0\] ram\[29\]\[0\] ram\[30\]\[0\] ram\[31\]\[0\] _0638_ _0628_
+ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1779_ _0575_ _0578_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__and2_1
X_3518_ clknet_leaf_9_clk _0080_ VGND VGND VPWR VPWR ram\[14\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3449_ _1723_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2820_ _1075_ ram\[35\]\[1\] _1377_ VGND VGND VPWR VPWR _1379_ sky130_fd_sc_hd__mux2_1
X_2751_ _1077_ net167 _1338_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2682_ _1300_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3303_ _1537_ net232 _1646_ VGND VGND VPWR VPWR _1647_ sky130_fd_sc_hd__mux2_1
X_3234_ _1451_ _1591_ VGND VGND VPWR VPWR _1610_ sky130_fd_sc_hd__nand2_4
X_3165_ _1537_ net194 _1572_ VGND VGND VPWR VPWR _1573_ sky130_fd_sc_hd__mux2_1
X_2116_ _0908_ _0909_ _0910_ _0644_ _0645_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__o221a_1
X_3096_ _1532_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__clkbuf_1
X_2047_ _0840_ _0841_ _0842_ _0595_ _0596_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__o221a_1
XFILLER_0_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2949_ _1395_ net354 _1452_ VGND VGND VPWR VPWR _1453_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold440 addr_reg\[0\] VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 ram\[46\]\[4\] VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 ram\[8\]\[1\] VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 ram\[49\]\[3\] VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 ram\[35\]\[0\] VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 ram\[45\]\[0\] VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_0_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3921_ clknet_leaf_38_clk _0477_ VGND VGND VPWR VPWR ram\[6\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_3852_ clknet_leaf_33_clk _0414_ VGND VGND VPWR VPWR ram\[56\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2803_ _1369_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_14_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3783_ clknet_leaf_21_clk _0345_ VGND VGND VPWR VPWR ram\[47\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2734_ _1077_ net143 _1329_ VGND VGND VPWR VPWR _1332_ sky130_fd_sc_hd__mux2_1
X_2665_ _1291_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__clkbuf_1
X_2596_ _1254_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3217_ _1441_ _1591_ VGND VGND VPWR VPWR _1601_ sky130_fd_sc_hd__nand2_4
XFILLER_0_66_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3148_ _1537_ net225 _1563_ VGND VGND VPWR VPWR _1564_ sky130_fd_sc_hd__mux2_1
X_3079_ _1523_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_59_Left_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_68_Left_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold270 ram\[1\]\[3\] VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 ram\[41\]\[2\] VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 ram\[54\]\[6\] VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_56_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2450_ _1170_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__clkbuf_1
X_2381_ _1077_ net528 _1128_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__mux2_1
Xinput5 addr[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_4
X_3002_ _1481_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3904_ clknet_leaf_28_clk _0466_ VGND VGND VPWR VPWR ram\[62\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3835_ clknet_leaf_28_clk _0397_ VGND VGND VPWR VPWR ram\[54\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3766_ clknet_leaf_20_clk _0328_ VGND VGND VPWR VPWR ram\[45\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2717_ net11 VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__buf_4
X_3697_ clknet_leaf_15_clk _0259_ VGND VGND VPWR VPWR ram\[36\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2648_ _1282_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__clkbuf_1
X_2579_ _1245_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1950_ _0618_ _0747_ _0621_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__o21a_1
X_1881_ _0675_ _0679_ _0598_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3620_ clknet_leaf_0_clk _0182_ VGND VGND VPWR VPWR ram\[27\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3551_ clknet_leaf_44_clk _0113_ VGND VGND VPWR VPWR ram\[18\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2502_ _1204_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3482_ clknet_leaf_10_clk _0044_ VGND VGND VPWR VPWR ram\[10\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2433_ _1160_ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__clkbuf_8
X_2364_ net309 _1062_ _1115_ VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2295_ net9 VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_67_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_10 _1323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3818_ clknet_leaf_29_clk _0380_ VGND VGND VPWR VPWR ram\[52\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_3749_ clknet_leaf_19_clk _0311_ VGND VGND VPWR VPWR ram\[43\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2080_ _0637_ _0871_ _0875_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_64_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2982_ _1051_ _1137_ VGND VGND VPWR VPWR _1470_ sky130_fd_sc_hd__nor2_4
XFILLER_0_56_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1933_ _0588_ ram\[48\]\[2\] VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3603_ clknet_leaf_1_clk _0165_ VGND VGND VPWR VPWR ram\[25\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_1864_ ram\[42\]\[1\] ram\[43\]\[1\] _0561_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__mux2_1
X_1795_ _0559_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__clkbuf_4
X_3534_ clknet_leaf_43_clk _0096_ VGND VGND VPWR VPWR ram\[16\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3465_ clknet_leaf_3_clk _0027_ VGND VGND VPWR VPWR ram\[29\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2416_ _1151_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__clkbuf_1
X_3396_ _1062_ net416 _1691_ VGND VGND VPWR VPWR _1696_ sky130_fd_sc_hd__mux2_1
X_2347_ net275 _1064_ _1104_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2278_ net253 _1064_ _1054_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3250_ _1618_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__clkbuf_1
X_3181_ _1498_ _1509_ VGND VGND VPWR VPWR _1581_ sky130_fd_sc_hd__nand2_4
X_2201_ _0934_ _0993_ _0621_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_77_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2132_ _0641_ ram\[9\]\[5\] _0652_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__a21o_1
X_2063_ ram\[20\]\[4\] ram\[21\]\[4\] _0629_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_22_Left_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2965_ _1127_ _1431_ VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__nand2_4
X_2896_ net412 _1315_ _1421_ VGND VGND VPWR VPWR _1423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1916_ ram\[44\]\[2\] ram\[45\]\[2\] ram\[46\]\[2\] ram\[47\]\[2\] _0548_ _0551_
+ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__mux4_1
X_1847_ _0637_ _0639_ _0646_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_31_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3517_ clknet_leaf_10_clk _0079_ VGND VGND VPWR VPWR ram\[14\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_1778_ ram\[32\]\[0\] ram\[33\]\[0\] ram\[34\]\[0\] ram\[35\]\[0\] _0576_ _0577_
+ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__mux4_1
X_3448_ _0540_ net24 net15 VGND VGND VPWR VPWR _1723_ sky130_fd_sc_hd__mux2_1
X_3379_ _1062_ net193 _1682_ VGND VGND VPWR VPWR _1687_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_40_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2750_ _1340_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2681_ _1083_ net427 _1294_ VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3302_ _1161_ _1591_ VGND VGND VPWR VPWR _1646_ sky130_fd_sc_hd__nand2_4
X_3233_ _1609_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__clkbuf_1
X_3164_ _1161_ _1509_ VGND VGND VPWR VPWR _1572_ sky130_fd_sc_hd__nand2_4
X_2115_ ram\[18\]\[5\] ram\[19\]\[5\] _0654_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__mux2_1
X_3095_ _1402_ ram\[50\]\[3\] _1528_ VGND VGND VPWR VPWR _1532_ sky130_fd_sc_hd__mux2_1
X_2046_ ram\[50\]\[4\] ram\[51\]\[4\] _0733_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2948_ _1451_ _1431_ VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__nand2_4
X_2879_ _1398_ net453 _1412_ VGND VGND VPWR VPWR _1414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold430 ram\[38\]\[1\] VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold463 ram\[27\]\[3\] VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 ram\[21\]\[1\] VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 ram\[44\]\[0\] VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 ram\[55\]\[6\] VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 ram\[43\]\[4\] VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 ram\[44\]\[4\] VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_0_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3920_ clknet_leaf_39_clk _0476_ VGND VGND VPWR VPWR ram\[6\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3851_ clknet_leaf_36_clk _0413_ VGND VGND VPWR VPWR ram\[56\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_3782_ clknet_leaf_20_clk _0344_ VGND VGND VPWR VPWR ram\[47\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2802_ net270 _1315_ _1367_ VGND VGND VPWR VPWR _1369_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2733_ _1331_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2664_ net198 _1194_ _1285_ VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__mux2_1
X_2595_ _1083_ net248 _1248_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3216_ _1600_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__clkbuf_1
X_3147_ _1149_ _1509_ VGND VGND VPWR VPWR _1563_ sky130_fd_sc_hd__nand2_4
X_3078_ net350 _1319_ _1519_ VGND VGND VPWR VPWR _1523_ sky130_fd_sc_hd__mux2_1
X_2029_ ram\[40\]\[4\] ram\[41\]\[4\] _0556_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold260 ram\[5\]\[4\] VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 ram\[54\]\[7\] VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 ram\[38\]\[0\] VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 ram\[21\]\[2\] VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_56_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2380_ _1130_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__clkbuf_1
Xinput6 addr[5] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
X_3001_ _1395_ net518 _1480_ VGND VGND VPWR VPWR _1481_ sky130_fd_sc_hd__mux2_1
X_3903_ clknet_leaf_32_clk _0465_ VGND VGND VPWR VPWR ram\[62\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_3834_ clknet_leaf_29_clk _0396_ VGND VGND VPWR VPWR ram\[54\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_62_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3765_ clknet_leaf_20_clk _0327_ VGND VGND VPWR VPWR ram\[45\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2716_ _1320_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__clkbuf_1
X_3696_ clknet_leaf_14_clk _0258_ VGND VGND VPWR VPWR ram\[36\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2647_ net347 _1194_ _1276_ VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2578_ _1083_ net351 _1239_ VGND VGND VPWR VPWR _1245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1880_ _0676_ _0677_ _0678_ _0595_ _0596_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__o221a_1
XFILLER_0_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3550_ clknet_leaf_43_clk _0112_ VGND VGND VPWR VPWR ram\[18\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2501_ net176 _1186_ _1202_ VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__mux2_1
X_3481_ clknet_leaf_36_clk _0043_ VGND VGND VPWR VPWR ram\[0\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2432_ net15 _1159_ VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2363_ _1119_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__clkbuf_1
X_2294_ _1076_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_67_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_11 _1406_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3817_ clknet_leaf_23_clk _0379_ VGND VGND VPWR VPWR ram\[51\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3748_ clknet_leaf_19_clk _0310_ VGND VGND VPWR VPWR ram\[43\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3679_ clknet_leaf_12_clk _0241_ VGND VGND VPWR VPWR ram\[34\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2981_ _1469_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_41_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_2
X_1932_ _0545_ _0729_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1863_ _0554_ _0661_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__or2_1
X_3602_ clknet_leaf_2_clk _0164_ VGND VGND VPWR VPWR ram\[25\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_1794_ ram\[50\]\[0\] ram\[51\]\[0\] _0593_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__mux2_1
X_3533_ clknet_leaf_42_clk _0095_ VGND VGND VPWR VPWR ram\[16\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3464_ clknet_leaf_2_clk _0026_ VGND VGND VPWR VPWR ram\[29\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2415_ _1070_ net241 _1150_ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__mux2_1
X_3395_ _1695_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2346_ _1109_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__clkbuf_1
X_2277_ net12 VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_32_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_74_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2200_ ram\[30\]\[7\] ram\[31\]\[7\] _0654_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3180_ _1580_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_77_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2131_ _0604_ ram\[8\]\[5\] VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__and2b_1
X_2062_ _0854_ _0856_ _0857_ _0626_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2964_ _1460_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_32_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1915_ _0673_ _0688_ _0713_ _0659_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_14_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_2
X_2895_ _1422_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1846_ _0640_ _0642_ _0643_ _0644_ _0645_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__o221a_1
X_1777_ _0549_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__buf_4
XFILLER_0_12_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3516_ clknet_leaf_9_clk _0078_ VGND VGND VPWR VPWR ram\[14\]\[2\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3447_ _1722_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__clkbuf_1
X_3378_ _1686_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__clkbuf_1
X_2329_ _1100_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2680_ _1299_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3301_ _1645_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__clkbuf_1
X_3232_ _1552_ net334 _1601_ VGND VGND VPWR VPWR _1609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_3_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_2
X_3163_ _1571_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__clkbuf_1
X_2114_ _0651_ ram\[17\]\[5\] _0652_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__a21o_1
X_3094_ _1531_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__clkbuf_1
X_2045_ _0568_ ram\[49\]\[4\] _0591_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2947_ _1051_ _1113_ VGND VGND VPWR VPWR _1451_ sky130_fd_sc_hd__nor2_4
X_2878_ _1413_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold420 ram\[31\]\[5\] VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__dlygate4sd3_1
X_1829_ _0000_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__buf_4
Xhold431 ram\[52\]\[5\] VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 addr_reg\[2\] VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold442 ram\[53\]\[7\] VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 ram\[27\]\[2\] VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 ram\[27\]\[4\] VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 ram\[47\]\[4\] VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold497 ram\[43\]\[0\] VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3850_ clknet_leaf_36_clk _0412_ VGND VGND VPWR VPWR ram\[56\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_3781_ clknet_leaf_20_clk _0343_ VGND VGND VPWR VPWR ram\[47\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2801_ _1368_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_14_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2732_ _1075_ net448 _1329_ VGND VGND VPWR VPWR _1331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2663_ _1290_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__clkbuf_1
X_2594_ _1253_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3215_ net108 _1327_ _1592_ VGND VGND VPWR VPWR _1600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3146_ _1562_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__clkbuf_1
X_3077_ _1522_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2028_ ram\[44\]\[4\] ram\[45\]\[4\] ram\[46\]\[4\] ram\[47\]\[4\] _0548_ _0551_
+ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__mux4_1
XFILLER_0_9_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold250 ram\[42\]\[2\] VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 ram\[34\]\[2\] VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold283 ram\[59\]\[3\] VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 ram\[51\]\[0\] VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 ram\[32\]\[3\] VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput7 data[0] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_4
XFILLER_0_36_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3000_ _1149_ _1431_ VGND VGND VPWR VPWR _1480_ sky130_fd_sc_hd__nand2_4
X_3902_ clknet_leaf_32_clk _0464_ VGND VGND VPWR VPWR ram\[62\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3833_ clknet_leaf_29_clk _0395_ VGND VGND VPWR VPWR ram\[53\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3764_ clknet_leaf_20_clk _0326_ VGND VGND VPWR VPWR ram\[45\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2715_ net114 _1319_ _1313_ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__mux2_1
X_3695_ clknet_leaf_15_clk _0257_ VGND VGND VPWR VPWR ram\[36\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2646_ _1281_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2577_ _1244_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3129_ _1553_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_53_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2500_ _1203_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__clkbuf_1
X_3480_ clknet_leaf_36_clk _0042_ VGND VGND VPWR VPWR ram\[0\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2431_ _0530_ net2 net3 VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__and3b_1
X_2362_ net313 _1060_ _1115_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__mux2_1
X_2293_ _1075_ net209 _1073_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_12 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3816_ clknet_leaf_23_clk _0378_ VGND VGND VPWR VPWR ram\[51\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3747_ clknet_leaf_19_clk _0309_ VGND VGND VPWR VPWR ram\[43\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_3678_ clknet_leaf_11_clk _0240_ VGND VGND VPWR VPWR ram\[34\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2629_ _1272_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2980_ _1410_ net189 _1461_ VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__mux2_1
X_1931_ ram\[52\]\[2\] ram\[53\]\[2\] ram\[54\]\[2\] ram\[55\]\[2\] _0547_ _0728_
+ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_72_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1862_ ram\[40\]\[1\] ram\[41\]\[1\] _0556_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput10 data[3] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_4
X_3601_ clknet_leaf_37_clk _0163_ VGND VGND VPWR VPWR ram\[24\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1793_ _0555_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__buf_4
X_3532_ clknet_leaf_42_clk _0094_ VGND VGND VPWR VPWR ram\[16\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3463_ clknet_leaf_1_clk _0025_ VGND VGND VPWR VPWR ram\[29\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2414_ _1125_ _1149_ VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__nand2_4
X_3394_ _1060_ net496 _1691_ VGND VGND VPWR VPWR _1695_ sky130_fd_sc_hd__mux2_1
X_2345_ net263 _1062_ _1104_ VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__mux2_1
X_2276_ _1063_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2130_ ram\[12\]\[5\] ram\[13\]\[5\] ram\[14\]\[5\] ram\[15\]\[5\] _0638_ _0624_
+ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__mux4_1
X_2061_ ram\[0\]\[4\] ram\[1\]\[4\] ram\[2\]\[4\] ram\[3\]\[4\] _0623_ _0634_ VGND
+ VGND VPWR VPWR _0857_ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2963_ _1410_ net78 _1452_ VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1914_ _0694_ _0700_ _0706_ _0712_ _0004_ _0543_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__mux4_2
XFILLER_0_44_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2894_ net77 _1312_ _1421_ VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1845_ _0563_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__buf_4
X_1776_ _0000_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__buf_4
XFILLER_0_71_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3515_ clknet_leaf_9_clk _0077_ VGND VGND VPWR VPWR ram\[14\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_3446_ net5 net282 net15 VGND VGND VPWR VPWR _1722_ sky130_fd_sc_hd__mux2_1
X_3377_ _1060_ net306 _1682_ VGND VGND VPWR VPWR _1686_ sky130_fd_sc_hd__mux2_1
X_2328_ net236 _1062_ _1095_ VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2259_ net15 VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__inv_4
XFILLER_0_47_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3300_ _1552_ net455 _1637_ VGND VGND VPWR VPWR _1645_ sky130_fd_sc_hd__mux2_1
X_3231_ _1608_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__clkbuf_1
X_3162_ _1552_ net465 _1563_ VGND VGND VPWR VPWR _1571_ sky130_fd_sc_hd__mux2_1
X_2113_ _0649_ ram\[16\]\[5\] VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__and2b_1
X_3093_ _1400_ ram\[50\]\[2\] _1528_ VGND VGND VPWR VPWR _1531_ sky130_fd_sc_hd__mux2_1
X_2044_ _0588_ ram\[48\]\[4\] VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__and2b_1
X_2946_ _1450_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__clkbuf_1
X_2877_ _1395_ net316 _1412_ VGND VGND VPWR VPWR _1413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1828_ _0549_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__buf_2
XFILLER_0_4_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold410 ram\[34\]\[0\] VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 ram\[27\]\[0\] VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__dlygate4sd3_1
X_1759_ _0001_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__inv_2
Xhold432 ram\[61\]\[7\] VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 ram\[37\]\[4\] VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold421 ram\[46\]\[2\] VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold465 ram\[0\]\[6\] VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 ram\[51\]\[6\] VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 ram\[47\]\[2\] VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 ram\[51\]\[2\] VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__dlygate4sd3_1
X_3429_ _1713_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_0_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3780_ clknet_leaf_20_clk _0342_ VGND VGND VPWR VPWR ram\[47\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2800_ net433 _1312_ _1367_ VGND VGND VPWR VPWR _1368_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2731_ _1330_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2662_ net153 _1192_ _1285_ VGND VGND VPWR VPWR _1290_ sky130_fd_sc_hd__mux2_1
X_2593_ _1081_ net165 _1248_ VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3214_ _1599_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_19_Left_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3145_ _1552_ net429 _1554_ VGND VGND VPWR VPWR _1562_ sky130_fd_sc_hd__mux2_1
X_3076_ net151 _1317_ _1519_ VGND VGND VPWR VPWR _1522_ sky130_fd_sc_hd__mux2_1
X_2027_ _0783_ _0798_ _0823_ _0659_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__a22o_1
XFILLER_0_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_28_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2929_ _1051_ _1200_ VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__nor2_4
XFILLER_0_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold240 ram\[0\]\[4\] VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 ram\[30\]\[3\] VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 ram\[33\]\[0\] VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 ram\[18\]\[0\] VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 ram\[19\]\[2\] VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 ram\[36\]\[2\] VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 data[1] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_19_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3901_ clknet_leaf_32_clk _0463_ VGND VGND VPWR VPWR ram\[62\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3832_ clknet_leaf_29_clk _0394_ VGND VGND VPWR VPWR ram\[53\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3763_ clknet_leaf_19_clk _0325_ VGND VGND VPWR VPWR ram\[45\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2714_ net10 VGND VGND VPWR VPWR _1319_ sky130_fd_sc_hd__buf_4
XFILLER_0_54_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3694_ clknet_leaf_16_clk _0256_ VGND VGND VPWR VPWR ram\[36\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2645_ net468 _1192_ _1276_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__mux2_1
X_2576_ _1081_ net199 _1239_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__mux2_1
X_3128_ _1552_ net524 _1538_ VGND VGND VPWR VPWR _1553_ sky130_fd_sc_hd__mux2_1
X_3059_ net422 _1317_ _1510_ VGND VGND VPWR VPWR _1513_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2430_ _1158_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__clkbuf_1
X_2361_ _1118_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2292_ net8 VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_67_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_13 _0585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3815_ clknet_leaf_28_clk _0377_ VGND VGND VPWR VPWR ram\[51\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3746_ clknet_leaf_19_clk _0308_ VGND VGND VPWR VPWR ram\[43\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3677_ clknet_leaf_11_clk _0239_ VGND VGND VPWR VPWR ram\[34\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2628_ net174 _1192_ _1267_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__mux2_1
X_2559_ _1234_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_38_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1930_ _0001_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_72_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1861_ ram\[44\]\[1\] ram\[45\]\[1\] ram\[46\]\[1\] ram\[47\]\[1\] _0548_ _0551_
+ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__mux4_1
Xinput11 data[4] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_4
X_3600_ clknet_leaf_38_clk _0162_ VGND VGND VPWR VPWR ram\[24\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3531_ clknet_leaf_44_clk _0093_ VGND VGND VPWR VPWR ram\[16\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1792_ _0590_ ram\[49\]\[0\] _0591_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3462_ clknet_leaf_7_clk _0024_ VGND VGND VPWR VPWR ram\[29\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3393_ _1694_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__clkbuf_1
X_2413_ _1148_ VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2344_ _1108_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__clkbuf_1
X_2275_ net331 _1062_ _1054_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3729_ clknet_leaf_15_clk _0291_ VGND VGND VPWR VPWR ram\[40\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2060_ _0618_ _0855_ _0621_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2962_ _1459_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_32_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1913_ _0637_ _0707_ _0711_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2893_ _0535_ _1053_ _0530_ _0533_ VGND VGND VPWR VPWR _1421_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1844_ _0559_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1775_ _0563_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3514_ clknet_leaf_8_clk _0076_ VGND VGND VPWR VPWR ram\[14\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_3445_ _1721_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__clkbuf_1
X_3376_ _1685_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__clkbuf_1
X_2327_ _1099_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2258_ _1049_ VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__inv_2
X_2189_ _0561_ ram\[36\]\[6\] VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3230_ _1550_ net35 _1601_ VGND VGND VPWR VPWR _1608_ sky130_fd_sc_hd__mux2_1
X_3161_ _1570_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__clkbuf_1
X_2112_ ram\[20\]\[5\] ram\[21\]\[5\] ram\[22\]\[5\] ram\[23\]\[5\] _0638_ _0628_
+ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__mux4_1
X_3092_ _1530_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__clkbuf_1
X_2043_ _0545_ _0838_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_45_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2945_ _1410_ net32 _1442_ VGND VGND VPWR VPWR _1450_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2876_ _1161_ _1376_ VGND VGND VPWR VPWR _1412_ sky130_fd_sc_hd__nand2_4
X_1827_ _0617_ _0622_ _0625_ _0626_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold400 ram\[58\]\[0\] VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold411 ram\[32\]\[7\] VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 ram\[57\]\[1\] VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold422 ram\[35\]\[6\] VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__dlygate4sd3_1
X_1758_ _0554_ _0557_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__or2_1
Xhold433 ram\[42\]\[3\] VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 ram\[18\]\[3\] VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 ram\[60\]\[1\] VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 ram\[37\]\[7\] VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold488 ram\[51\]\[4\] VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__dlygate4sd3_1
X_3428_ net286 net10 _1709_ VGND VGND VPWR VPWR _1713_ sky130_fd_sc_hd__mux2_1
Xhold499 ram\[11\]\[0\] VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__dlygate4sd3_1
X_3359_ _1676_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_13_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2730_ _1070_ net266 _1329_ VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2661_ _1289_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__clkbuf_1
X_2592_ _1252_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3213_ net367 _1325_ _1592_ VGND VGND VPWR VPWR _1599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3144_ _1561_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__clkbuf_1
X_3075_ _1521_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__clkbuf_1
X_2026_ _0804_ _0810_ _0816_ _0822_ _0004_ _0611_ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__mux4_2
XFILLER_0_9_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2928_ _1440_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2859_ _1400_ net104 _1396_ VGND VGND VPWR VPWR _1401_ sky130_fd_sc_hd__mux2_1
Xhold230 ram\[7\]\[5\] VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 ram\[0\]\[5\] VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 ram\[9\]\[7\] VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 ram\[15\]\[5\] VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 ram\[40\]\[4\] VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 ram\[39\]\[3\] VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 ram\[10\]\[2\] VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 data[2] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_19_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3900_ clknet_leaf_32_clk _0462_ VGND VGND VPWR VPWR ram\[62\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3831_ clknet_leaf_30_clk _0393_ VGND VGND VPWR VPWR ram\[53\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_3762_ clknet_leaf_20_clk _0324_ VGND VGND VPWR VPWR ram\[45\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2713_ _1318_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__clkbuf_1
X_3693_ clknet_leaf_16_clk _0255_ VGND VGND VPWR VPWR ram\[36\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2644_ _1280_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__clkbuf_1
X_2575_ _1243_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3127_ net14 VGND VGND VPWR VPWR _1552_ sky130_fd_sc_hd__buf_2
X_3058_ _1512_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2009_ _0628_ _0805_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_53_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_47_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2360_ net297 _1058_ _1115_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2291_ _1074_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Left_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_44_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_14 _0600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3814_ clknet_leaf_30_clk _0376_ VGND VGND VPWR VPWR ram\[51\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3745_ clknet_leaf_21_clk _0307_ VGND VGND VPWR VPWR ram\[42\]\[7\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_65_Left_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3676_ clknet_leaf_11_clk _0238_ VGND VGND VPWR VPWR ram\[34\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2627_ _1271_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2558_ net84 _1192_ _1229_ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2489_ _1195_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_74_Left_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_35_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_21_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_26_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_56_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1860_ _0582_ _0613_ _0658_ _0659_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__a22o_1
Xinput12 data[5] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_4
X_1791_ _0549_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3530_ clknet_leaf_43_clk _0092_ VGND VGND VPWR VPWR ram\[16\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3461_ clknet_leaf_7_clk _0023_ VGND VGND VPWR VPWR ram\[29\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_3392_ _1058_ net529 _1691_ VGND VGND VPWR VPWR _1694_ sky130_fd_sc_hd__mux2_1
X_2412_ net15 _1072_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__and2_1
X_2343_ net65 _1060_ _1104_ VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__mux2_1
X_2274_ net11 VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__buf_4
XFILLER_0_74_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_17_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_35_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1989_ _0588_ ram\[48\]\[3\] VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__and2b_1
XFILLER_0_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3728_ clknet_leaf_24_clk _0290_ VGND VGND VPWR VPWR ram\[40\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3659_ clknet_leaf_17_clk _0221_ VGND VGND VPWR VPWR ram\[32\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2961_ _1408_ net333 _1452_ VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1912_ _0708_ _0709_ _0710_ _0644_ _0645_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__o221a_1
XFILLER_0_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2892_ _1420_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1843_ ram\[10\]\[0\] ram\[11\]\[0\] _0576_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1774_ _0569_ _0571_ _0572_ _0560_ _0573_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3513_ clknet_leaf_13_clk _0075_ VGND VGND VPWR VPWR ram\[13\]\[7\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_6_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_2
X_3444_ _0537_ net197 _0531_ VGND VGND VPWR VPWR _1721_ sky130_fd_sc_hd__mux2_1
X_3375_ _1058_ net290 _1682_ VGND VGND VPWR VPWR _1685_ sky130_fd_sc_hd__mux2_1
X_2326_ net52 _1060_ _1095_ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__mux2_1
X_2257_ _0530_ _0533_ _0535_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__and3_2
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2188_ _0977_ _0981_ _0542_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3160_ _1550_ net461 _1563_ VGND VGND VPWR VPWR _1570_ sky130_fd_sc_hd__mux2_1
X_2111_ _0584_ _0898_ _0905_ _0005_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__o31a_1
Xhold1 addr_reg\[5\] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dlygate4sd3_1
X_3091_ _1398_ ram\[50\]\[1\] _1528_ VGND VGND VPWR VPWR _1530_ sky130_fd_sc_hd__mux2_1
X_2042_ ram\[52\]\[4\] ram\[53\]\[4\] ram\[54\]\[4\] ram\[55\]\[4\] _0547_ _0728_
+ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2944_ _1449_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2875_ _1411_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1826_ _0563_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold401 ram\[61\]\[2\] VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold423 ram\[43\]\[2\] VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 ram\[25\]\[4\] VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 ram\[11\]\[6\] VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 ram\[13\]\[3\] VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__dlygate4sd3_1
X_1757_ ram\[40\]\[0\] ram\[41\]\[0\] _0556_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__mux2_1
Xhold456 ram\[57\]\[0\] VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 ram\[45\]\[2\] VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 ram\[11\]\[3\] VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold489 ram\[45\]\[6\] VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__dlygate4sd3_1
X_3427_ _1712_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__clkbuf_1
X_3358_ _1058_ net124 _1673_ VGND VGND VPWR VPWR _1676_ sky130_fd_sc_hd__mux2_1
X_2309_ _1086_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__clkbuf_1
X_3289_ _1639_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_0_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2660_ net149 _1190_ _1285_ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2591_ _1079_ net211 _1248_ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3212_ _1598_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3143_ _1550_ net358 _1554_ VGND VGND VPWR VPWR _1561_ sky130_fd_sc_hd__mux2_1
X_3074_ net74 _1315_ _1519_ VGND VGND VPWR VPWR _1521_ sky130_fd_sc_hd__mux2_1
X_2025_ _0637_ _0817_ _0821_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2927_ net152 _1327_ _1432_ VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2858_ net9 VGND VGND VPWR VPWR _1400_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1809_ ram\[56\]\[0\] ram\[57\]\[0\] ram\[58\]\[0\] ram\[59\]\[0\] _0608_ _0553_
+ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__mux4_1
Xhold220 ram\[9\]\[6\] VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__dlygate4sd3_1
X_2789_ net187 _1319_ _1358_ VGND VGND VPWR VPWR _1362_ sky130_fd_sc_hd__mux2_1
Xhold253 ram\[16\]\[1\] VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 ram\[52\]\[1\] VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 ram\[30\]\[4\] VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 ram\[5\]\[3\] VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 ram\[23\]\[6\] VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 ram\[10\]\[4\] VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 ram\[46\]\[7\] VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_56_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3830_ clknet_leaf_31_clk _0392_ VGND VGND VPWR VPWR ram\[53\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3761_ clknet_leaf_22_clk _0323_ VGND VGND VPWR VPWR ram\[44\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2712_ net117 _1317_ _1313_ VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__mux2_1
X_3692_ clknet_leaf_16_clk _0254_ VGND VGND VPWR VPWR ram\[36\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2643_ net426 _1190_ _1276_ VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__mux2_1
X_2574_ _1079_ net106 _1239_ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__mux2_1
X_3126_ _1551_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__clkbuf_1
X_3057_ net105 _1315_ _1510_ VGND VGND VPWR VPWR _1512_ sky130_fd_sc_hd__mux2_1
X_2008_ ram\[20\]\[3\] ram\[21\]\[3\] _0629_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3959_ clknet_leaf_38_clk _0515_ VGND VGND VPWR VPWR ram\[19\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_61_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2290_ _1070_ net484 _1073_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3813_ clknet_leaf_28_clk _0375_ VGND VGND VPWR VPWR ram\[51\]\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_15 _1064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3744_ clknet_leaf_23_clk _0306_ VGND VGND VPWR VPWR ram\[42\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3675_ clknet_leaf_11_clk _0237_ VGND VGND VPWR VPWR ram\[34\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2626_ net381 _1190_ _1267_ VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2557_ _1233_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2488_ net186 _1194_ _1184_ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__mux2_1
X_3109_ net8 VGND VGND VPWR VPWR _1540_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_66_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput13 data[6] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_4
X_1790_ _0567_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__buf_4
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3460_ clknet_leaf_6_clk _0022_ VGND VGND VPWR VPWR ram\[29\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3391_ _1693_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__clkbuf_1
X_2411_ _1147_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__clkbuf_1
X_2342_ _1107_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__clkbuf_1
X_2273_ _1061_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1988_ _0545_ _0784_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__and2_1
X_3727_ clknet_leaf_15_clk _0289_ VGND VGND VPWR VPWR ram\[40\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3658_ clknet_leaf_16_clk _0220_ VGND VGND VPWR VPWR ram\[32\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2609_ _1261_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__clkbuf_1
X_3589_ clknet_leaf_5_clk _0151_ VGND VGND VPWR VPWR ram\[23\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_26_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2960_ _1458_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1911_ ram\[26\]\[1\] ram\[27\]\[1\] _0619_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__mux2_1
X_2891_ _1410_ net389 _1412_ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1842_ _0641_ ram\[9\]\[0\] _0550_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1773_ _0544_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__buf_4
XFILLER_0_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3512_ clknet_leaf_13_clk _0074_ VGND VGND VPWR VPWR ram\[13\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3443_ _1720_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__clkbuf_1
X_3374_ _1684_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__clkbuf_1
X_2325_ _1098_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__clkbuf_1
X_2256_ net7 VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__buf_4
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2187_ _0978_ _0979_ _0980_ _0934_ _0944_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_48_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2110_ _0902_ _0904_ _0542_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__o21a_1
X_3090_ _1529_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__clkbuf_1
Xhold2 ram\[40\]\[6\] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2041_ _0543_ _0829_ _0836_ _0581_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_45_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2943_ _1408_ net99 _1442_ VGND VGND VPWR VPWR _1449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2874_ _1410_ net500 _1396_ VGND VGND VPWR VPWR _1411_ sky130_fd_sc_hd__mux2_1
X_1825_ ram\[0\]\[0\] ram\[1\]\[0\] ram\[2\]\[0\] ram\[3\]\[0\] _0623_ _0624_ VGND
+ VGND VPWR VPWR _0625_ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold402 ram\[18\]\[5\] VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1756_ _0555_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__buf_4
Xhold435 ram\[63\]\[3\] VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold413 ram\[5\]\[6\] VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold424 ram\[49\]\[0\] VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 ram\[58\]\[1\] VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 ram\[52\]\[3\] VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 ram\[42\]\[4\] VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3426_ net344 net9 _1709_ VGND VGND VPWR VPWR _1712_ sky130_fd_sc_hd__mux2_1
Xhold479 ram\[35\]\[4\] VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__dlygate4sd3_1
X_3357_ _1675_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__clkbuf_1
X_2308_ _1085_ net404 _1073_ VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__mux2_1
X_3288_ _1540_ ram\[61\]\[1\] _1637_ VGND VGND VPWR VPWR _1639_ sky130_fd_sc_hd__mux2_1
X_2239_ _0543_ _1024_ _1031_ _0584_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__a211o_1
XFILLER_0_45_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2590_ _1251_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3211_ net86 _1323_ _1592_ VGND VGND VPWR VPWR _1598_ sky130_fd_sc_hd__mux2_1
X_3142_ _1560_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__clkbuf_1
X_3073_ _1520_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__clkbuf_1
X_2024_ _0818_ _0819_ _0820_ _0644_ _0645_ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__o221a_1
X_2926_ _1439_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2857_ _1399_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__clkbuf_1
X_1808_ _0000_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__clkbuf_8
X_2788_ _1361_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__clkbuf_1
Xhold210 ram\[62\]\[3\] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold221 ram\[24\]\[1\] VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 ram\[61\]\[6\] VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__dlygate4sd3_1
X_1739_ net6 VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__buf_2
Xhold243 ram\[30\]\[0\] VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 ram\[40\]\[2\] VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 ram\[39\]\[5\] VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 ram\[13\]\[4\] VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 ram\[10\]\[1\] VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__dlygate4sd3_1
X_3409_ _1058_ net296 _1700_ VGND VGND VPWR VPWR _1703_ sky130_fd_sc_hd__mux2_1
Xhold298 ram\[47\]\[1\] VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3760_ clknet_leaf_22_clk _0322_ VGND VGND VPWR VPWR ram\[44\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2711_ net9 VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__buf_4
XFILLER_0_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3691_ clknet_leaf_17_clk _0253_ VGND VGND VPWR VPWR ram\[36\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2642_ _1279_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2573_ _1242_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3125_ _1550_ net499 _1538_ VGND VGND VPWR VPWR _1551_ sky130_fd_sc_hd__mux2_1
X_3056_ _1511_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2007_ _0800_ _0802_ _0803_ _0626_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3958_ clknet_leaf_39_clk _0514_ VGND VGND VPWR VPWR ram\[19\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_61_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2909_ _1429_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__clkbuf_1
X_3889_ clknet_leaf_28_clk _0451_ VGND VGND VPWR VPWR ram\[60\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3812_ clknet_leaf_30_clk _0374_ VGND VGND VPWR VPWR ram\[51\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_16 _1315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3743_ clknet_leaf_21_clk _0305_ VGND VGND VPWR VPWR ram\[42\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3674_ clknet_leaf_11_clk _0236_ VGND VGND VPWR VPWR ram\[34\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2625_ _1270_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2556_ net130 _1190_ _1229_ VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__mux2_1
X_2487_ net12 VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__buf_2
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3108_ _1539_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_66_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3039_ _1501_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_38_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput14 data[7] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2410_ net384 _1068_ _1139_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__mux2_1
X_3390_ _1056_ net400 _1691_ VGND VGND VPWR VPWR _1693_ sky130_fd_sc_hd__mux2_1
X_2341_ net146 _1058_ _1104_ VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__mux2_1
X_2272_ net289 _1060_ _1054_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1987_ ram\[52\]\[3\] ram\[53\]\[3\] ram\[54\]\[3\] ram\[55\]\[3\] _0547_ _0728_
+ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__mux4_1
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3726_ clknet_leaf_15_clk _0288_ VGND VGND VPWR VPWR ram\[40\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3657_ clknet_leaf_3_clk _0219_ VGND VGND VPWR VPWR ram\[31\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3588_ clknet_leaf_4_clk _0150_ VGND VGND VPWR VPWR ram\[23\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2608_ net100 _1190_ _1257_ VGND VGND VPWR VPWR _1261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2539_ net293 _1190_ _1220_ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1910_ _0651_ ram\[25\]\[1\] _0652_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__a21o_1
X_2890_ _1419_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_32_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1841_ _0555_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1772_ ram\[38\]\[0\] ram\[39\]\[0\] _0556_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3511_ clknet_leaf_8_clk _0073_ VGND VGND VPWR VPWR ram\[13\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_3442_ _0535_ net476 _0531_ VGND VGND VPWR VPWR _1720_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3373_ _1056_ net397 _1682_ VGND VGND VPWR VPWR _1684_ sky130_fd_sc_hd__mux2_1
X_2324_ net390 _1058_ _1095_ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__mux2_1
X_2255_ _0659_ _1004_ _1018_ _1032_ _1047_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__a32o_1
XFILLER_0_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2186_ ram\[42\]\[6\] ram\[43\]\[6\] _0733_ VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3709_ clknet_leaf_18_clk _0271_ VGND VGND VPWR VPWR ram\[38\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3 ram\[41\]\[3\] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dlygate4sd3_1
X_2040_ _0833_ _0835_ _0598_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_29_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2942_ _1448_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2873_ net14 VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__buf_2
X_1824_ _0549_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__buf_4
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1755_ _0000_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__clkbuf_4
Xhold436 ram\[61\]\[3\] VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold403 ram\[25\]\[3\] VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 ram\[30\]\[1\] VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 ram\[14\]\[5\] VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 ram\[60\]\[4\] VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold458 ram\[45\]\[3\] VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold447 ram\[45\]\[1\] VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3425_ _1711_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__clkbuf_1
X_3356_ _1056_ net494 _1673_ VGND VGND VPWR VPWR _1675_ sky130_fd_sc_hd__mux2_1
X_3287_ _1638_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__clkbuf_1
X_2307_ net13 VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__buf_2
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2238_ _1028_ _1030_ _0598_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__o21ba_1
X_2169_ ram\[56\]\[6\] ram\[57\]\[6\] _0593_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3210_ _1597_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__clkbuf_1
X_3141_ _1548_ net454 _1554_ VGND VGND VPWR VPWR _1560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3072_ net258 _1312_ _1519_ VGND VGND VPWR VPWR _1520_ sky130_fd_sc_hd__mux2_1
X_2023_ ram\[26\]\[3\] ram\[27\]\[3\] _0619_ VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__mux2_1
X_2925_ net25 _1325_ _1432_ VGND VGND VPWR VPWR _1439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2856_ _1398_ net517 _1396_ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__mux2_1
X_1807_ _0601_ _0603_ _0605_ _0606_ _0573_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_13_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2787_ net349 _1317_ _1358_ VGND VGND VPWR VPWR _1361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold211 ram\[62\]\[5\] VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold200 ram\[53\]\[4\] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 ram\[4\]\[7\] VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 ram\[28\]\[1\] VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1738_ _0539_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__clkbuf_1
Xhold222 ram\[35\]\[5\] VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 ram\[60\]\[3\] VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 ram\[7\]\[3\] VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold255 ram\[58\]\[7\] VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3408_ _1702_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__clkbuf_1
Xhold288 ram\[20\]\[5\] VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 ram\[8\]\[7\] VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__dlygate4sd3_1
X_3339_ net44 net8 _1664_ VGND VGND VPWR VPWR _1666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2710_ _1316_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3690_ clknet_leaf_16_clk _0252_ VGND VGND VPWR VPWR ram\[36\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_10_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2641_ net365 _1188_ _1276_ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__mux2_1
X_2572_ _1077_ net305 _1239_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3124_ net13 VGND VGND VPWR VPWR _1550_ sky130_fd_sc_hd__buf_2
X_3055_ net406 _1312_ _1510_ VGND VGND VPWR VPWR _1511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2006_ ram\[0\]\[3\] ram\[1\]\[3\] ram\[2\]\[3\] ram\[3\]\[3\] _0623_ _0634_ VGND
+ VGND VPWR VPWR _0803_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_53_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3957_ clknet_leaf_43_clk _0513_ VGND VGND VPWR VPWR ram\[19\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2908_ net220 _1327_ _1421_ VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3888_ clknet_leaf_28_clk _0450_ VGND VGND VPWR VPWR ram\[60\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2839_ net307 _1317_ _1386_ VGND VGND VPWR VPWR _1389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_38_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_16_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_25_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3811_ clknet_leaf_28_clk _0373_ VGND VGND VPWR VPWR ram\[51\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_17 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3742_ clknet_leaf_20_clk _0304_ VGND VGND VPWR VPWR ram\[42\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3673_ clknet_leaf_15_clk _0235_ VGND VGND VPWR VPWR ram\[33\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2624_ net513 _1188_ _1267_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_34_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2555_ _1232_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2486_ _1193_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__clkbuf_1
X_3107_ _1537_ net317 _1538_ VGND VGND VPWR VPWR _1539_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3038_ _1398_ net321 _1499_ VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_52_Left_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Left_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput15 we VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_70_Left_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2340_ _1106_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2271_ net10 VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_63_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1986_ _0543_ _0775_ _0782_ _0581_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__a211o_1
XFILLER_0_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3725_ clknet_leaf_17_clk _0287_ VGND VGND VPWR VPWR ram\[40\]\[3\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_9_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_2
X_3656_ clknet_leaf_3_clk _0218_ VGND VGND VPWR VPWR ram\[31\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3587_ clknet_leaf_2_clk _0149_ VGND VGND VPWR VPWR ram\[23\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2607_ _1260_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2538_ _1223_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__clkbuf_1
X_2469_ net7 VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1840_ _0604_ ram\[8\]\[0\] VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3510_ clknet_leaf_8_clk _0072_ VGND VGND VPWR VPWR ram\[13\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_1771_ _0548_ ram\[37\]\[0\] _0570_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__a21o_1
X_3441_ _1719_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__clkbuf_1
X_3372_ _1683_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__clkbuf_1
X_2323_ _1097_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__clkbuf_1
X_2254_ _0581_ _1039_ _1046_ _0005_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__o31a_1
XFILLER_0_79_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2185_ _0600_ ram\[41\]\[6\] _0577_ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1969_ _0764_ _0765_ _0766_ _0644_ _0645_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__o221a_1
X_3708_ clknet_leaf_16_clk _0270_ VGND VGND VPWR VPWR ram\[38\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3639_ clknet_leaf_41_clk _0201_ VGND VGND VPWR VPWR ram\[2\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold4 ram\[41\]\[5\] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlygate4sd3_1
X_2941_ _1406_ net27 _1442_ VGND VGND VPWR VPWR _1448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2872_ _1409_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__clkbuf_1
X_1823_ _0567_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__buf_4
X_1754_ _0553_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__buf_2
XFILLER_0_20_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold426 ram\[27\]\[6\] VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold404 ram\[27\]\[5\] VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold415 ram\[62\]\[7\] VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 ram\[50\]\[7\] VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__dlygate4sd3_1
X_3424_ net388 net8 _1709_ VGND VGND VPWR VPWR _1711_ sky130_fd_sc_hd__mux2_1
Xhold459 ram\[44\]\[3\] VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 ram\[44\]\[1\] VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__dlygate4sd3_1
X_3355_ _1674_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3286_ _1537_ net531 _1637_ VGND VGND VPWR VPWR _1638_ sky130_fd_sc_hd__mux2_1
X_2306_ _1084_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__clkbuf_1
X_2237_ _0944_ _1029_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2168_ ram\[60\]\[6\] ram\[61\]\[6\] ram\[62\]\[6\] ram\[63\]\[6\] _0548_ _0551_
+ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_0_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2099_ _0588_ ram\[48\]\[5\] VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3140_ _1559_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_8_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3071_ _1053_ _1137_ VGND VGND VPWR VPWR _1519_ sky130_fd_sc_hd__nor2_4
X_2022_ _0651_ ram\[25\]\[3\] _0652_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3973_ clknet_leaf_26_clk _0529_ VGND VGND VPWR VPWR addr_reg\[5\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2924_ _1438_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__clkbuf_1
X_2855_ net8 VGND VGND VPWR VPWR _1398_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1806_ _0559_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2786_ _1360_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__clkbuf_1
Xhold201 ram\[12\]\[6\] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold223 ram\[4\]\[4\] VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 ram\[3\]\[4\] VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 ram\[62\]\[4\] VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__dlygate4sd3_1
X_1737_ net5 net282 _0531_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__mux2_1
Xhold267 ram\[59\]\[2\] VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 ram\[4\]\[6\] VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 ram\[24\]\[7\] VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 ram\[30\]\[7\] VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3407_ _1056_ net374 _1700_ VGND VGND VPWR VPWR _1702_ sky130_fd_sc_hd__mux2_1
Xhold289 ram\[7\]\[7\] VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__dlygate4sd3_1
X_3338_ _1665_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3269_ _1537_ net451 _1628_ VGND VGND VPWR VPWR _1629_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2640_ _1278_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_10_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2571_ _1241_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3123_ _1549_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__clkbuf_1
X_3054_ _1094_ _1509_ VGND VGND VPWR VPWR _1510_ sky130_fd_sc_hd__nor2b_4
X_2005_ _0618_ _0801_ _0621_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_53_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3956_ clknet_leaf_43_clk _0512_ VGND VGND VPWR VPWR ram\[19\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2907_ _1428_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3887_ clknet_leaf_32_clk _0449_ VGND VGND VPWR VPWR ram\[60\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2838_ _1388_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__clkbuf_1
X_2769_ _1351_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3810_ clknet_leaf_28_clk _0372_ VGND VGND VPWR VPWR ram\[51\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_18 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3741_ clknet_leaf_19_clk _0303_ VGND VGND VPWR VPWR ram\[42\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3672_ clknet_leaf_14_clk _0234_ VGND VGND VPWR VPWR ram\[33\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2623_ _1269_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2554_ net49 _1188_ _1229_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2485_ net217 _1192_ _1184_ VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__mux2_1
X_3106_ _1127_ _1509_ VGND VGND VPWR VPWR _1538_ sky130_fd_sc_hd__nand2_4
XFILLER_0_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3037_ _1500_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3939_ clknet_leaf_34_clk _0495_ VGND VGND VPWR VPWR ram\[59\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2270_ _1059_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_63_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1985_ _0779_ _0781_ _0598_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__o21ba_1
X_3724_ clknet_leaf_17_clk _0286_ VGND VGND VPWR VPWR ram\[40\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3655_ clknet_leaf_8_clk _0217_ VGND VGND VPWR VPWR ram\[31\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2606_ net67 _1188_ _1257_ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__mux2_1
X_3586_ clknet_leaf_4_clk _0148_ VGND VGND VPWR VPWR ram\[23\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2537_ net136 _1188_ _1220_ VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2468_ _1180_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2399_ _1141_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1770_ _0549_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3440_ _0533_ net385 _0531_ VGND VGND VPWR VPWR _1719_ sky130_fd_sc_hd__mux2_1
X_3371_ _1048_ net188 _1682_ VGND VGND VPWR VPWR _1683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2322_ net474 _1056_ _1095_ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2253_ _1043_ _1045_ _0003_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_18_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2184_ _0651_ ram\[40\]\[6\] VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_48_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1968_ ram\[26\]\[2\] ram\[27\]\[2\] _0619_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3707_ clknet_leaf_17_clk _0269_ VGND VGND VPWR VPWR ram\[38\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_1899_ _0618_ _0697_ _0544_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__o21a_1
X_3638_ clknet_leaf_41_clk _0200_ VGND VGND VPWR VPWR ram\[2\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3569_ clknet_leaf_3_clk _0131_ VGND VGND VPWR VPWR ram\[20\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold5 ram\[58\]\[6\] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2940_ _1447_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__clkbuf_1
X_2871_ _1408_ net48 _1396_ VGND VGND VPWR VPWR _1409_ sky130_fd_sc_hd__mux2_1
X_1822_ _0618_ _0620_ _0621_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1753_ _0549_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__buf_4
XFILLER_0_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold416 ram\[61\]\[4\] VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold427 ram\[52\]\[0\] VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold405 ram\[45\]\[4\] VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 ram\[53\]\[6\] VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 ram\[35\]\[7\] VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__dlygate4sd3_1
X_3423_ _1710_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__clkbuf_1
X_3354_ _1048_ net76 _1673_ VGND VGND VPWR VPWR _1674_ sky130_fd_sc_hd__mux2_1
X_2305_ _1083_ net407 _1073_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__mux2_1
X_3285_ _1149_ _1591_ VGND VGND VPWR VPWR _1637_ sky130_fd_sc_hd__nand2_4
X_2236_ ram\[48\]\[7\] ram\[49\]\[7\] ram\[50\]\[7\] ram\[51\]\[7\] _0629_ _0652_
+ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2167_ _0611_ _0953_ _0960_ _0581_ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_0_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2098_ _0545_ _0892_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3070_ _1518_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__clkbuf_1
X_2021_ _0649_ ram\[24\]\[3\] VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__and2b_1
XFILLER_0_49_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3972_ clknet_leaf_14_clk _0528_ VGND VGND VPWR VPWR addr_reg\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2923_ net207 _1323_ _1432_ VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2854_ _1397_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2785_ net116 _1315_ _1358_ VGND VGND VPWR VPWR _1360_ sky130_fd_sc_hd__mux2_1
X_1805_ ram\[62\]\[0\] ram\[63\]\[0\] _0604_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold202 ram\[53\]\[0\] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__dlygate4sd3_1
X_1736_ _0538_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__clkbuf_1
Xhold235 ram\[4\]\[0\] VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 ram\[47\]\[7\] VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 ram\[8\]\[4\] VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold246 ram\[54\]\[1\] VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 ram\[31\]\[7\] VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 ram\[38\]\[4\] VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__dlygate4sd3_1
X_3406_ _1701_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__clkbuf_1
Xhold279 ram\[55\]\[1\] VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3337_ net175 net7 _1664_ VGND VGND VPWR VPWR _1665_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _1470_ _1591_ VGND VGND VPWR VPWR _1628_ sky130_fd_sc_hd__nand2_4
X_2219_ _0623_ ram\[5\]\[7\] _0577_ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__a21o_1
X_3199_ _1590_ VGND VGND VPWR VPWR _1591_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_56_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2570_ _1075_ net464 _1239_ VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3122_ _1548_ net356 _1538_ VGND VGND VPWR VPWR _1549_ sky130_fd_sc_hd__mux2_1
X_3053_ _1508_ VGND VGND VPWR VPWR _1509_ sky130_fd_sc_hd__buf_6
X_2004_ ram\[6\]\[3\] ram\[7\]\[3\] _0619_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3955_ clknet_leaf_42_clk _0511_ VGND VGND VPWR VPWR ram\[19\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2906_ net164 _1325_ _1421_ VGND VGND VPWR VPWR _1428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3886_ clknet_leaf_32_clk _0448_ VGND VGND VPWR VPWR ram\[60\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2837_ net112 _1315_ _1386_ VGND VGND VPWR VPWR _1388_ sky130_fd_sc_hd__mux2_1
X_2768_ net249 _1315_ _1349_ VGND VGND VPWR VPWR _1351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2699_ _1309_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_69_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3740_ clknet_leaf_19_clk _0302_ VGND VGND VPWR VPWR ram\[42\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3671_ clknet_leaf_12_clk _0233_ VGND VGND VPWR VPWR ram\[33\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2622_ net244 _1186_ _1267_ VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__mux2_1
X_2553_ _1231_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__clkbuf_1
X_2484_ net11 VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3105_ net7 VGND VGND VPWR VPWR _1537_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_66_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3036_ _1395_ net516 _1499_ VGND VGND VPWR VPWR _1500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3938_ clknet_leaf_35_clk _0494_ VGND VGND VPWR VPWR ram\[59\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3869_ clknet_leaf_34_clk _0431_ VGND VGND VPWR VPWR ram\[58\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1984_ _0575_ _0780_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_71_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3723_ clknet_leaf_17_clk _0285_ VGND VGND VPWR VPWR ram\[40\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_3654_ clknet_leaf_7_clk _0216_ VGND VGND VPWR VPWR ram\[31\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2605_ _1259_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__clkbuf_1
X_3585_ clknet_leaf_4_clk _0147_ VGND VGND VPWR VPWR ram\[22\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2536_ _1222_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__clkbuf_1
X_2467_ net221 _1068_ _1172_ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2398_ net42 _1056_ _1139_ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3019_ _1490_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_77_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3370_ _1127_ _1591_ VGND VGND VPWR VPWR _1682_ sky130_fd_sc_hd__nand2_4
X_2321_ _1096_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__clkbuf_1
X_2252_ _0944_ _1044_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2183_ _0545_ _0976_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_48_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1967_ _0651_ ram\[25\]\[2\] _0652_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__a21o_1
X_3706_ clknet_leaf_17_clk _0268_ VGND VGND VPWR VPWR ram\[38\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_1898_ ram\[22\]\[1\] ram\[23\]\[1\] _0608_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__mux2_1
X_3637_ clknet_leaf_40_clk _0199_ VGND VGND VPWR VPWR ram\[2\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3568_ clknet_leaf_3_clk _0130_ VGND VGND VPWR VPWR ram\[20\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2519_ _1213_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__clkbuf_1
X_3499_ clknet_leaf_9_clk _0061_ VGND VGND VPWR VPWR ram\[12\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Left_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_58_Left_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold6 ram\[1\]\[0\] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2870_ net13 VGND VGND VPWR VPWR _1408_ sky130_fd_sc_hd__buf_2
X_1821_ _0544_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_2
X_1752_ ram\[44\]\[0\] ram\[45\]\[0\] ram\[46\]\[0\] ram\[47\]\[0\] _0548_ _0551_
+ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__mux4_1
XFILLER_0_25_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold406 ram\[52\]\[7\] VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 ram\[43\]\[1\] VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold428 ram\[60\]\[0\] VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3422_ net401 net7 _1709_ VGND VGND VPWR VPWR _1710_ sky130_fd_sc_hd__mux2_1
Xhold439 ram\[12\]\[3\] VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3353_ _1498_ _1591_ VGND VGND VPWR VPWR _1673_ sky130_fd_sc_hd__nand2_4
XFILLER_0_29_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3284_ _1636_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__clkbuf_1
X_2304_ net12 VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__buf_2
X_2235_ _1025_ _1026_ _1027_ _0595_ _0585_ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__o221a_1
X_2166_ _0957_ _0959_ _0003_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_0_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2097_ ram\[52\]\[5\] ram\[53\]\[5\] ram\[54\]\[5\] ram\[55\]\[5\] _0547_ _0728_
+ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2999_ _1479_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2020_ ram\[28\]\[3\] ram\[29\]\[3\] ram\[30\]\[3\] ram\[31\]\[3\] _0638_ _0624_
+ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__mux4_1
X_3971_ clknet_leaf_14_clk _0527_ VGND VGND VPWR VPWR addr_reg\[3\] sky130_fd_sc_hd__dfxtp_1
X_2922_ _1437_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2853_ _1395_ ram\[37\]\[0\] _1396_ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1804_ _0555_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__buf_4
X_2784_ _1359_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__clkbuf_1
X_1735_ _0537_ net197 _0531_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__mux2_1
Xhold214 ram\[0\]\[7\] VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold203 ram\[26\]\[7\] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 ram\[22\]\[5\] VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 ram\[19\]\[4\] VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 ram\[22\]\[1\] VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 ram\[31\]\[1\] VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 ram\[34\]\[1\] VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__dlygate4sd3_1
X_3405_ _1048_ net441 _1700_ VGND VGND VPWR VPWR _1701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3336_ _1053_ _1159_ VGND VGND VPWR VPWR _1664_ sky130_fd_sc_hd__nor2b_4
X_3267_ _1627_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2218_ _0641_ ram\[4\]\[7\] VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__and2b_1
X_3198_ _0537_ net5 net6 VGND VGND VPWR VPWR _1590_ sky130_fd_sc_hd__and3_1
X_2149_ ram\[18\]\[6\] ram\[19\]\[6\] _0654_ VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3121_ net12 VGND VGND VPWR VPWR _1548_ sky130_fd_sc_hd__buf_2
X_3052_ _1089_ net5 net6 VGND VGND VPWR VPWR _1508_ sky130_fd_sc_hd__and3_1
X_2003_ _0614_ _0799_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_18_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3954_ clknet_leaf_43_clk _0510_ VGND VGND VPWR VPWR ram\[19\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3885_ clknet_leaf_32_clk _0447_ VGND VGND VPWR VPWR ram\[60\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2905_ _1427_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_61_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2836_ _1387_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2767_ _1350_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__clkbuf_1
X_2698_ net409 _1194_ _1303_ VGND VGND VPWR VPWR _1309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3319_ _1091_ _1201_ VGND VGND VPWR VPWR _1655_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_69_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3670_ clknet_leaf_11_clk _0232_ VGND VGND VPWR VPWR ram\[33\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2621_ _1268_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2552_ net338 _1186_ _1229_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__mux2_1
X_2483_ _1191_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3104_ _1536_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__clkbuf_1
X_3035_ _1498_ _1431_ VGND VGND VPWR VPWR _1499_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_66_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3937_ clknet_leaf_36_clk _0493_ VGND VGND VPWR VPWR ram\[59\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_3868_ clknet_leaf_35_clk _0430_ VGND VGND VPWR VPWR ram\[58\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3799_ clknet_leaf_35_clk _0361_ VGND VGND VPWR VPWR ram\[4\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2819_ _1378_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1983_ ram\[32\]\[3\] ram\[33\]\[3\] ram\[34\]\[3\] ram\[35\]\[3\] _0576_ _0577_
+ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__mux4_1
X_3722_ clknet_leaf_17_clk _0284_ VGND VGND VPWR VPWR ram\[40\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_3653_ clknet_leaf_7_clk _0215_ VGND VGND VPWR VPWR ram\[31\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2604_ net190 _1186_ _1257_ VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__mux2_1
X_3584_ clknet_leaf_3_clk _0146_ VGND VGND VPWR VPWR ram\[22\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2535_ net222 _1186_ _1220_ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2466_ _1179_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__clkbuf_1
X_2397_ _1140_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3018_ _1395_ net505 _1489_ VGND VGND VPWR VPWR _1490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2320_ net170 _1048_ _1095_ VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__mux2_1
X_2251_ ram\[32\]\[7\] ram\[33\]\[7\] ram\[34\]\[7\] ram\[35\]\[7\] _0629_ _0550_
+ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__mux4_1
XFILLER_0_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2182_ ram\[44\]\[6\] ram\[45\]\[6\] ram\[46\]\[6\] ram\[47\]\[6\] _0567_ _0728_
+ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1966_ _0649_ ram\[24\]\[2\] VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3705_ clknet_leaf_23_clk _0267_ VGND VGND VPWR VPWR ram\[37\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_1897_ _0628_ _0695_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__or2_1
X_3636_ clknet_leaf_42_clk _0198_ VGND VGND VPWR VPWR ram\[2\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3567_ clknet_leaf_1_clk _0129_ VGND VGND VPWR VPWR ram\[20\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2518_ net410 _1186_ _1211_ VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3498_ clknet_leaf_8_clk _0060_ VGND VGND VPWR VPWR ram\[12\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2449_ _1087_ net421 _1162_ VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold7 ram\[56\]\[2\] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_45_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1820_ ram\[6\]\[0\] ram\[7\]\[0\] _0619_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1751_ _0550_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__buf_4
Xhold418 ram\[19\]\[0\] VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold407 ram\[14\]\[3\] VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__dlygate4sd3_1
X_3421_ _1171_ _1348_ VGND VGND VPWR VPWR _1709_ sky130_fd_sc_hd__nor2_4
Xhold429 ram\[36\]\[3\] VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3352_ _1672_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2303_ _1082_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__clkbuf_1
X_3283_ _1552_ net379 _1628_ VGND VGND VPWR VPWR _1636_ sky130_fd_sc_hd__mux2_1
X_2234_ ram\[54\]\[7\] ram\[55\]\[7\] _0593_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__mux2_1
X_2165_ _0645_ _0958_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__and2_1
X_2096_ _0543_ _0883_ _0890_ _0581_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2998_ _1410_ net185 _1471_ VGND VGND VPWR VPWR _1479_ sky130_fd_sc_hd__mux2_1
X_1949_ ram\[6\]\[2\] ram\[7\]\[2\] _0619_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3619_ clknet_leaf_0_clk _0181_ VGND VGND VPWR VPWR ram\[27\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_8_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3970_ clknet_leaf_37_clk _0526_ VGND VGND VPWR VPWR addr_reg\[2\] sky130_fd_sc_hd__dfxtp_1
X_2921_ net308 _1321_ _1432_ VGND VGND VPWR VPWR _1437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2852_ _1149_ _1376_ VGND VGND VPWR VPWR _1396_ sky130_fd_sc_hd__nand2_4
XFILLER_0_72_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1803_ _0602_ ram\[61\]\[0\] _0570_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_13_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2783_ net274 _1312_ _1358_ VGND VGND VPWR VPWR _1359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1734_ net4 VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__buf_2
Xhold226 ram\[32\]\[1\] VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold204 ram\[5\]\[2\] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 ram\[15\]\[0\] VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 ram\[26\]\[6\] VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__dlygate4sd3_1
X_3404_ _1127_ _1238_ VGND VGND VPWR VPWR _1700_ sky130_fd_sc_hd__nand2_4
Xhold259 addr_reg\[4\] VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 ram\[37\]\[5\] VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3335_ _1663_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__clkbuf_1
X_3266_ net420 net14 _1619_ VGND VGND VPWR VPWR _1627_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2217_ _0546_ _1005_ _1007_ _1009_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3197_ _1589_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_77_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2148_ _0588_ ram\[17\]\[6\] _0553_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__a21o_1
X_2079_ _0872_ _0873_ _0874_ _0644_ _0645_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__o221a_1
XFILLER_0_48_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3120_ _1547_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__clkbuf_1
X_3051_ _1507_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__clkbuf_1
X_2002_ ram\[4\]\[3\] ram\[5\]\[3\] _0615_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3953_ clknet_leaf_44_clk _0509_ VGND VGND VPWR VPWR ram\[19\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3884_ clknet_leaf_31_clk _0446_ VGND VGND VPWR VPWR ram\[60\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2904_ net192 _1323_ _1421_ VGND VGND VPWR VPWR _1427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2835_ net183 _1312_ _1386_ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2766_ net179 _1312_ _1349_ VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2697_ _1308_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3318_ _1654_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__clkbuf_1
X_3249_ _1552_ net278 _1610_ VGND VGND VPWR VPWR _1618_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2620_ net145 _1181_ _1267_ VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2551_ _1230_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2482_ net110 _1190_ _1184_ VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__mux2_1
X_3103_ _1410_ net460 _1528_ VGND VGND VPWR VPWR _1536_ sky130_fd_sc_hd__mux2_1
X_3034_ _1051_ _1050_ VGND VGND VPWR VPWR _1498_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_66_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3936_ clknet_leaf_35_clk _0492_ VGND VGND VPWR VPWR ram\[59\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_3867_ clknet_leaf_36_clk _0429_ VGND VGND VPWR VPWR ram\[58\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_3798_ clknet_leaf_40_clk _0360_ VGND VGND VPWR VPWR ram\[4\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2818_ _1070_ net507 _1377_ VGND VGND VPWR VPWR _1378_ sky130_fd_sc_hd__mux2_1
X_2749_ _1075_ net292 _1338_ VGND VGND VPWR VPWR _1340_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1982_ _0776_ _0777_ _0778_ _0606_ _0573_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_71_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3721_ clknet_leaf_37_clk _0283_ VGND VGND VPWR VPWR ram\[3\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3652_ clknet_leaf_7_clk _0214_ VGND VGND VPWR VPWR ram\[31\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3583_ clknet_leaf_1_clk _0145_ VGND VGND VPWR VPWR ram\[22\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2603_ _1258_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__clkbuf_1
X_2534_ _1221_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2465_ net31 _1066_ _1172_ VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__mux2_1
X_2396_ net262 _1048_ _1139_ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3017_ _1161_ _1431_ VGND VGND VPWR VPWR _1489_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_34_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3919_ clknet_leaf_13_clk _0475_ VGND VGND VPWR VPWR ram\[9\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2250_ _1040_ _1041_ _1042_ _0934_ _0585_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__o221a_1
X_2181_ _0543_ _0967_ _0974_ _0584_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_48_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1965_ ram\[28\]\[2\] ram\[29\]\[2\] ram\[30\]\[2\] ram\[31\]\[2\] _0638_ _0628_
+ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__mux4_1
XFILLER_0_28_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3704_ clknet_leaf_24_clk _0266_ VGND VGND VPWR VPWR ram\[37\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_1896_ ram\[20\]\[1\] ram\[21\]\[1\] _0629_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__mux2_1
X_3635_ clknet_leaf_42_clk _0197_ VGND VGND VPWR VPWR ram\[2\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3566_ clknet_leaf_6_clk _0128_ VGND VGND VPWR VPWR ram\[20\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2517_ _1212_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__clkbuf_1
X_3497_ clknet_leaf_12_clk _0059_ VGND VGND VPWR VPWR ram\[11\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2448_ _1169_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_39_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2379_ _1075_ net473 _1128_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold8 ram\[15\]\[6\] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_73_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1750_ _0549_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__buf_4
XFILLER_0_25_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold408 ram\[54\]\[5\] VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__dlygate4sd3_1
X_3420_ _1708_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__clkbuf_1
Xhold419 ram\[55\]\[3\] VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3351_ net208 net14 _1664_ VGND VGND VPWR VPWR _1672_ sky130_fd_sc_hd__mux2_1
X_2302_ _1081_ net119 _1073_ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__mux2_1
X_3282_ _1635_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__clkbuf_1
X_2233_ _0590_ ram\[53\]\[7\] _0591_ VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__a21o_1
X_2164_ ram\[0\]\[6\] ram\[1\]\[6\] ram\[2\]\[6\] ram\[3\]\[6\] _0547_ _0728_ VGND
+ VGND VPWR VPWR _0958_ sky130_fd_sc_hd__mux4_1
X_2095_ _0887_ _0889_ _0598_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_48_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2997_ _1478_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__clkbuf_1
X_1948_ _0614_ _0745_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1879_ ram\[50\]\[1\] ram\[51\]\[1\] _0593_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3618_ clknet_leaf_1_clk _0180_ VGND VGND VPWR VPWR ram\[27\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3549_ clknet_leaf_43_clk _0111_ VGND VGND VPWR VPWR ram\[18\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_58_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2920_ _1436_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2851_ net7 VGND VGND VPWR VPWR _1395_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1802_ _0547_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__buf_4
X_2782_ _1201_ _1348_ VGND VGND VPWR VPWR _1358_ sky130_fd_sc_hd__nor2_4
X_1733_ _0536_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold205 ram\[57\]\[4\] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold216 ram\[33\]\[7\] VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 ram\[58\]\[2\] VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 ram\[48\]\[4\] VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 ram\[26\]\[2\] VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__dlygate4sd3_1
X_3403_ _1699_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3334_ net264 net14 _1655_ VGND VGND VPWR VPWR _1663_ sky130_fd_sc_hd__mux2_1
X_3265_ _1626_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__clkbuf_1
X_2216_ _0595_ _1008_ _0944_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__o21a_1
X_3196_ _1552_ net372 _1581_ VGND VGND VPWR VPWR _1589_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2147_ _0641_ ram\[16\]\[6\] VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__and2b_1
X_2078_ ram\[26\]\[4\] ram\[27\]\[4\] _0619_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_12_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3050_ _1410_ net247 _1499_ VGND VGND VPWR VPWR _1507_ sky130_fd_sc_hd__mux2_1
X_2001_ _0584_ _0790_ _0797_ _0005_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_18_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3952_ clknet_leaf_43_clk _0508_ VGND VGND VPWR VPWR ram\[19\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2903_ _1426_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__clkbuf_1
X_3883_ clknet_leaf_30_clk _0445_ VGND VGND VPWR VPWR ram\[60\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2834_ _1138_ _1348_ VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__nor2_4
X_2765_ _1094_ _1348_ VGND VGND VPWR VPWR _1349_ sky130_fd_sc_hd__nor2_4
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2696_ net75 _1192_ _1303_ VGND VGND VPWR VPWR _1308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3317_ _1552_ net438 _1646_ VGND VGND VPWR VPWR _1654_ sky130_fd_sc_hd__mux2_1
X_3248_ _1617_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_69_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3179_ _1552_ net294 _1572_ VGND VGND VPWR VPWR _1580_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_443 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2550_ net88 _1181_ _1229_ VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__mux2_1
X_2481_ net10 VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3102_ _1535_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__clkbuf_1
X_3033_ _1497_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_66_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3935_ clknet_leaf_28_clk _0491_ VGND VGND VPWR VPWR ram\[63\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3866_ clknet_leaf_35_clk _0428_ VGND VGND VPWR VPWR ram\[58\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3797_ clknet_leaf_40_clk _0359_ VGND VGND VPWR VPWR ram\[4\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2817_ _1127_ _1376_ VGND VGND VPWR VPWR _1377_ sky130_fd_sc_hd__nand2_4
XFILLER_0_5_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2748_ _1339_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__clkbuf_1
X_2679_ _1081_ net487 _1294_ VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3720_ clknet_leaf_35_clk _0282_ VGND VGND VPWR VPWR ram\[3\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_1981_ ram\[38\]\[3\] ram\[39\]\[3\] _0649_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_40_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_70_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3651_ clknet_leaf_0_clk _0213_ VGND VGND VPWR VPWR ram\[31\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2602_ net62 _1181_ _1257_ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__mux2_1
X_3582_ clknet_leaf_5_clk _0144_ VGND VGND VPWR VPWR ram\[22\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2533_ net29 _1181_ _1220_ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2464_ _1178_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2395_ _1091_ _1138_ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_79_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3016_ _1488_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_31_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_2
X_3918_ clknet_leaf_14_clk _0474_ VGND VGND VPWR VPWR ram\[9\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3849_ clknet_leaf_22_clk _0411_ VGND VGND VPWR VPWR ram\[55\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_22_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2180_ _0971_ _0973_ _0598_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_76_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_13_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_2
X_1964_ _0637_ _0757_ _0761_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3703_ clknet_leaf_21_clk _0265_ VGND VGND VPWR VPWR ram\[37\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_3634_ clknet_leaf_42_clk _0196_ VGND VGND VPWR VPWR ram\[2\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_1895_ _0690_ _0692_ _0693_ _0626_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__a22o_1
X_3565_ clknet_leaf_6_clk _0127_ VGND VGND VPWR VPWR ram\[20\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2516_ net318 _1181_ _1211_ VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__mux2_1
X_3496_ clknet_leaf_13_clk _0058_ VGND VGND VPWR VPWR ram\[11\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2447_ _1085_ net161 _1162_ VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2378_ _1129_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_39_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_18_Left_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold9 ram\[41\]\[7\] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_2_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold409 ram\[54\]\[3\] VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3350_ _1671_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__clkbuf_1
X_2301_ net11 VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__clkbuf_4
X_3281_ _1550_ net403 _1628_ VGND VGND VPWR VPWR _1635_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_2_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_2
X_2232_ _0623_ ram\[52\]\[7\] VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__and2b_1
X_2163_ _0954_ _0955_ _0956_ _0934_ _0545_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__o221a_1
XFILLER_0_45_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2094_ _0575_ _0888_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2996_ _1408_ net157 _1471_ VGND VGND VPWR VPWR _1478_ sky130_fd_sc_hd__mux2_1
X_1947_ ram\[4\]\[2\] ram\[5\]\[2\] _0615_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__mux2_1
X_1878_ _0590_ ram\[49\]\[1\] _0591_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3617_ clknet_leaf_2_clk _0179_ VGND VGND VPWR VPWR ram\[26\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3548_ clknet_leaf_43_clk _0110_ VGND VGND VPWR VPWR ram\[18\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3479_ clknet_leaf_40_clk _0041_ VGND VGND VPWR VPWR ram\[0\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2850_ _1394_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__clkbuf_1
X_1801_ _0600_ ram\[60\]\[0\] VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__and2b_1
XFILLER_0_72_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2781_ _1357_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1732_ _0535_ addr_reg\[2\] _0531_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__mux2_1
Xhold206 ram\[54\]\[4\] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 ram\[57\]\[2\] VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__dlygate4sd3_1
X_3402_ _1068_ net46 _1691_ VGND VGND VPWR VPWR _1699_ sky130_fd_sc_hd__mux2_1
Xhold228 ram\[13\]\[7\] VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 ram\[12\]\[0\] VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3333_ _1662_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3264_ net436 net13 _1619_ VGND VGND VPWR VPWR _1626_ sky130_fd_sc_hd__mux2_1
X_2215_ ram\[10\]\[7\] ram\[11\]\[7\] _0593_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__mux2_1
X_3195_ _1588_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2146_ _0621_ _0939_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__and2_1
X_2077_ _0651_ ram\[25\]\[4\] _0652_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2979_ _1468_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2000_ _0794_ _0796_ _0542_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_18_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3951_ clknet_leaf_25_clk _0507_ VGND VGND VPWR VPWR ram\[49\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2902_ net257 _1321_ _1421_ VGND VGND VPWR VPWR _1426_ sky130_fd_sc_hd__mux2_1
X_3882_ clknet_leaf_30_clk _0444_ VGND VGND VPWR VPWR ram\[60\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2833_ _1385_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__clkbuf_1
X_2764_ _1347_ VGND VGND VPWR VPWR _1348_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2695_ _1307_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__clkbuf_1
X_3316_ _1653_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3247_ _1550_ net28 _1610_ VGND VGND VPWR VPWR _1617_ sky130_fd_sc_hd__mux2_1
X_3178_ _1579_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__clkbuf_1
X_2129_ _0920_ _0922_ _0923_ _0626_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2480_ _1189_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3101_ _1408_ net493 _1528_ VGND VGND VPWR VPWR _1535_ sky130_fd_sc_hd__mux2_1
X_3032_ _1410_ net320 _1489_ VGND VGND VPWR VPWR _1497_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3934_ clknet_leaf_28_clk _0490_ VGND VGND VPWR VPWR ram\[63\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3865_ clknet_leaf_27_clk _0427_ VGND VGND VPWR VPWR ram\[57\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2816_ _1089_ _1124_ _0540_ VGND VGND VPWR VPWR _1376_ sky130_fd_sc_hd__and3_4
XFILLER_0_73_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3796_ clknet_leaf_35_clk _0358_ VGND VGND VPWR VPWR ram\[4\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2747_ _1070_ net355 _1338_ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2678_ _1298_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1980_ _0602_ ram\[37\]\[3\] _0570_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__a21o_1
X_3650_ clknet_leaf_8_clk _0212_ VGND VGND VPWR VPWR ram\[31\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2601_ _1171_ _1183_ VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__nor2_4
X_3581_ clknet_leaf_5_clk _0143_ VGND VGND VPWR VPWR ram\[22\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2532_ _1053_ _1200_ VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__nor2_4
X_2463_ net319 _1064_ _1172_ VGND VGND VPWR VPWR _1178_ sky130_fd_sc_hd__mux2_1
X_2394_ _1051_ _1137_ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__or2_4
XFILLER_0_48_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3015_ _1410_ net368 _1480_ VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3917_ clknet_leaf_4_clk _0473_ VGND VGND VPWR VPWR ram\[9\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_3848_ clknet_leaf_29_clk _0410_ VGND VGND VPWR VPWR ram\[55\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3779_ clknet_leaf_19_clk _0341_ VGND VGND VPWR VPWR ram\[47\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1963_ _0758_ _0759_ _0760_ _0644_ _0563_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__o221a_1
X_1894_ ram\[0\]\[1\] ram\[1\]\[1\] ram\[2\]\[1\] ram\[3\]\[1\] _0623_ _0624_ VGND
+ VGND VPWR VPWR _0693_ sky130_fd_sc_hd__mux4_1
XFILLER_0_55_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3702_ clknet_leaf_19_clk _0264_ VGND VGND VPWR VPWR ram\[37\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3633_ clknet_leaf_3_clk _0195_ VGND VGND VPWR VPWR ram\[28\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3564_ clknet_leaf_6_clk _0126_ VGND VGND VPWR VPWR ram\[20\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2515_ _1114_ _1183_ VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__nor2_4
X_3495_ clknet_leaf_5_clk _0057_ VGND VGND VPWR VPWR ram\[11\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2446_ _1168_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2377_ _1070_ net522 _1128_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3280_ _1634_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__clkbuf_1
X_2300_ _1080_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2231_ _0546_ _1019_ _1021_ _1023_ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__a22o_1
X_2162_ ram\[6\]\[6\] ram\[7\]\[6\] _0654_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__mux2_1
X_2093_ ram\[32\]\[5\] ram\[33\]\[5\] ram\[34\]\[5\] ram\[35\]\[5\] _0608_ _0553_
+ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2995_ _1477_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__clkbuf_1
X_1946_ _0584_ _0736_ _0743_ _0005_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__o31a_1
X_1877_ _0588_ ram\[48\]\[1\] VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3616_ clknet_leaf_2_clk _0178_ VGND VGND VPWR VPWR ram\[26\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3547_ clknet_leaf_44_clk _0109_ VGND VGND VPWR VPWR ram\[18\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_3478_ clknet_leaf_41_clk _0040_ VGND VGND VPWR VPWR ram\[0\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2429_ _1087_ net251 _1150_ VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1800_ _0567_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__buf_4
XFILLER_0_25_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2780_ net434 _1327_ _1349_ VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1731_ net3 VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__clkbuf_2
Xhold207 ram\[14\]\[4\] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__dlygate4sd3_1
X_3401_ _1698_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__clkbuf_1
Xhold229 ram\[43\]\[6\] VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 ram\[13\]\[0\] VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__dlygate4sd3_1
X_3332_ net243 net13 _1655_ VGND VGND VPWR VPWR _1662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3263_ _1625_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_37_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3194_ _1550_ net497 _1581_ VGND VGND VPWR VPWR _1588_ sky130_fd_sc_hd__mux2_1
X_2214_ _0554_ _1006_ VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__or2_1
X_2145_ ram\[20\]\[6\] ram\[21\]\[6\] ram\[22\]\[6\] ram\[23\]\[6\] _0567_ _0728_
+ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__mux4_1
X_2076_ _0649_ ram\[24\]\[4\] VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__and2b_1
XFILLER_0_72_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_46_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2978_ _1408_ net252 _1461_ VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1929_ _0543_ _0719_ _0726_ _0581_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__a211o_1
XFILLER_0_71_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_55_Left_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_64_Left_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Left_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold90 ram\[23\]\[4\] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dlygate4sd3_1
X_3950_ clknet_leaf_23_clk _0506_ VGND VGND VPWR VPWR ram\[49\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2901_ _1425_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__clkbuf_1
X_3881_ clknet_leaf_37_clk _0443_ VGND VGND VPWR VPWR ram\[5\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2832_ _1087_ net472 _1377_ VGND VGND VPWR VPWR _1385_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2763_ _0537_ net5 _0540_ VGND VGND VPWR VPWR _1347_ sky130_fd_sc_hd__or3b_1
XFILLER_0_53_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2694_ net66 _1190_ _1303_ VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3315_ _1550_ net411 _1646_ VGND VGND VPWR VPWR _1653_ sky130_fd_sc_hd__mux2_1
X_3246_ _1616_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3177_ _1550_ net315 _1572_ VGND VGND VPWR VPWR _1579_ sky130_fd_sc_hd__mux2_1
X_2128_ ram\[0\]\[5\] ram\[1\]\[5\] ram\[2\]\[5\] ram\[3\]\[5\] _0623_ _0634_ VGND
+ VGND VPWR VPWR _0923_ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2059_ ram\[6\]\[4\] ram\[7\]\[4\] _0619_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3100_ _1534_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__clkbuf_1
X_3031_ _1496_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_66_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3933_ clknet_leaf_33_clk _0489_ VGND VGND VPWR VPWR ram\[63\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_3864_ clknet_leaf_26_clk _0426_ VGND VGND VPWR VPWR ram\[57\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2815_ _1375_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__clkbuf_1
X_3795_ clknet_leaf_39_clk _0357_ VGND VGND VPWR VPWR ram\[4\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2746_ _1049_ _1071_ VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__nand2_4
X_2677_ _1079_ net486 _1294_ VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3229_ _1607_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold390 ram\[59\]\[5\] VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_63_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3580_ clknet_leaf_5_clk _0142_ VGND VGND VPWR VPWR ram\[22\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2600_ _1256_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__clkbuf_1
X_2531_ _1219_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2462_ _1177_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__clkbuf_1
X_2393_ _0530_ _0533_ _0535_ VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__or3b_4
X_3014_ _1487_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3916_ clknet_leaf_12_clk _0472_ VGND VGND VPWR VPWR ram\[9\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3847_ clknet_leaf_30_clk _0409_ VGND VGND VPWR VPWR ram\[55\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3778_ clknet_leaf_20_clk _0340_ VGND VGND VPWR VPWR ram\[47\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2729_ _1071_ _1159_ VGND VGND VPWR VPWR _1329_ sky130_fd_sc_hd__nand2_4
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1962_ ram\[10\]\[2\] ram\[11\]\[2\] _0576_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__mux2_1
X_1893_ _0618_ _0691_ _0621_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3701_ clknet_leaf_18_clk _0263_ VGND VGND VPWR VPWR ram\[37\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_3632_ clknet_leaf_2_clk _0194_ VGND VGND VPWR VPWR ram\[28\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3563_ clknet_leaf_1_clk _0125_ VGND VGND VPWR VPWR ram\[20\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2514_ _1210_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__clkbuf_1
X_3494_ clknet_leaf_10_clk _0056_ VGND VGND VPWR VPWR ram\[11\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2445_ _1083_ net437 _1162_ VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2376_ _1125_ _1127_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__nand2_4
XFILLER_0_78_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2230_ _0560_ _1022_ _0575_ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__o21a_1
X_2161_ _0623_ ram\[5\]\[6\] _0577_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2092_ _0884_ _0885_ _0886_ _0606_ _0573_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__o221a_1
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2994_ _1406_ net92 _1471_ VGND VGND VPWR VPWR _1477_ sky130_fd_sc_hd__mux2_1
X_1945_ _0740_ _0742_ _0542_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1876_ _0585_ _0674_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__and2_1
X_3615_ clknet_leaf_44_clk _0177_ VGND VGND VPWR VPWR ram\[26\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_3546_ clknet_leaf_43_clk _0108_ VGND VGND VPWR VPWR ram\[18\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3477_ clknet_leaf_34_clk _0039_ VGND VGND VPWR VPWR ram\[0\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2428_ _1157_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__clkbuf_1
X_2359_ _1117_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1730_ _0534_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold208 ram\[9\]\[2\] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3400_ _1066_ net483 _1691_ VGND VGND VPWR VPWR _1698_ sky130_fd_sc_hd__mux2_1
Xhold219 ram\[10\]\[6\] VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3331_ _1661_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__clkbuf_1
X_3262_ net182 net12 _1619_ VGND VGND VPWR VPWR _1625_ sky130_fd_sc_hd__mux2_1
X_3193_ _1587_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__clkbuf_1
X_2213_ ram\[8\]\[7\] ram\[9\]\[7\] _0733_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__mux2_1
X_2144_ _0933_ _0936_ _0937_ _0626_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__a22o_1
X_2075_ ram\[28\]\[4\] ram\[29\]\[4\] ram\[30\]\[4\] ram\[31\]\[4\] _0638_ _0624_
+ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__mux4_1
XFILLER_0_29_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2977_ _1467_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__clkbuf_1
X_1928_ _0723_ _0725_ _0542_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__o21ba_1
X_1859_ _0005_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__inv_2
X_3529_ clknet_leaf_13_clk _0091_ VGND VGND VPWR VPWR ram\[15\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold80 ram\[60\]\[2\] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 ram\[2\]\[3\] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dlygate4sd3_1
X_2900_ net214 _1319_ _1421_ VGND VGND VPWR VPWR _1425_ sky130_fd_sc_hd__mux2_1
X_3880_ clknet_leaf_36_clk _0442_ VGND VGND VPWR VPWR ram\[5\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2831_ _1384_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__clkbuf_1
X_2762_ _1346_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2693_ _1306_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__clkbuf_1
X_3314_ _1652_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__clkbuf_1
X_3245_ _1548_ net79 _1610_ VGND VGND VPWR VPWR _1616_ sky130_fd_sc_hd__mux2_1
X_3176_ _1578_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_16_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2127_ _0618_ _0921_ _0621_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2058_ _0614_ _0853_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_52_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3030_ _1408_ net402 _1489_ VGND VGND VPWR VPWR _1496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_43_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_2
X_3932_ clknet_leaf_34_clk _0488_ VGND VGND VPWR VPWR ram\[63\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3863_ clknet_leaf_33_clk _0425_ VGND VGND VPWR VPWR ram\[57\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2814_ net59 _1327_ _1367_ VGND VGND VPWR VPWR _1375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3794_ clknet_leaf_40_clk _0356_ VGND VGND VPWR VPWR ram\[4\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2745_ _1337_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2676_ _1297_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3228_ _1548_ net173 _1601_ VGND VGND VPWR VPWR _1607_ sky130_fd_sc_hd__mux2_1
X_3159_ _1569_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_29_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_34_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_76_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold380 ram\[60\]\[6\] VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 ram\[53\]\[5\] VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_63_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_67_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2530_ net41 _1198_ _1211_ VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2461_ net129 _1062_ _1172_ VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__mux2_1
X_2392_ _1136_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3013_ _1408_ net512 _1480_ VGND VGND VPWR VPWR _1487_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_16_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3915_ clknet_leaf_12_clk _0471_ VGND VGND VPWR VPWR ram\[9\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3846_ clknet_leaf_31_clk _0408_ VGND VGND VPWR VPWR ram\[55\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3777_ clknet_leaf_22_clk _0339_ VGND VGND VPWR VPWR ram\[46\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2728_ _1328_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__clkbuf_1
X_2659_ _1288_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1961_ _0641_ ram\[9\]\[2\] _0550_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__a21o_1
X_3700_ clknet_leaf_18_clk _0262_ VGND VGND VPWR VPWR ram\[37\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_1892_ ram\[6\]\[1\] ram\[7\]\[1\] _0619_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3631_ clknet_leaf_1_clk _0193_ VGND VGND VPWR VPWR ram\[28\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3562_ clknet_leaf_6_clk _0124_ VGND VGND VPWR VPWR ram\[20\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2513_ net90 _1198_ _1202_ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3493_ clknet_leaf_11_clk _0055_ VGND VGND VPWR VPWR ram\[11\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_2
X_2444_ _1167_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__clkbuf_1
X_2375_ _1126_ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3829_ clknet_leaf_29_clk _0391_ VGND VGND VPWR VPWR ram\[53\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2160_ _0641_ ram\[4\]\[6\] VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__and2b_1
X_2091_ ram\[38\]\[5\] ram\[39\]\[5\] _0649_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2993_ _1476_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__clkbuf_1
X_1944_ _0596_ _0741_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3614_ clknet_leaf_0_clk _0176_ VGND VGND VPWR VPWR ram\[26\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_1875_ ram\[52\]\[1\] ram\[53\]\[1\] ram\[54\]\[1\] ram\[55\]\[1\] _0547_ _0550_
+ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3545_ clknet_leaf_38_clk _0107_ VGND VGND VPWR VPWR ram\[17\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3476_ clknet_leaf_41_clk _0038_ VGND VGND VPWR VPWR ram\[0\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2427_ _1085_ net343 _1150_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2358_ net277 _1056_ _1115_ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__mux2_1
X_2289_ _1071_ _1072_ VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_50_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold209 ram\[62\]\[0\] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__dlygate4sd3_1
X_3330_ net89 net12 _1655_ VGND VGND VPWR VPWR _1661_ sky130_fd_sc_hd__mux2_1
X_3261_ _1624_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__clkbuf_1
X_3192_ _1548_ net417 _1581_ VGND VGND VPWR VPWR _1587_ sky130_fd_sc_hd__mux2_1
X_2212_ ram\[12\]\[7\] ram\[13\]\[7\] ram\[14\]\[7\] ram\[15\]\[7\] _0590_ _0614_
+ VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__mux4_1
X_2143_ ram\[24\]\[6\] ram\[25\]\[6\] ram\[26\]\[6\] ram\[27\]\[6\] _0602_ _0614_
+ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__mux4_1
X_2074_ _0573_ _0865_ _0869_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2976_ _1406_ net324 _1461_ VGND VGND VPWR VPWR _1467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1927_ _0575_ _0724_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1858_ _0627_ _0636_ _0647_ _0657_ _0004_ _0543_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__mux4_2
XFILLER_0_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1789_ _0588_ ram\[48\]\[0\] VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__and2b_1
X_3528_ clknet_leaf_4_clk _0090_ VGND VGND VPWR VPWR ram\[15\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3459_ clknet_leaf_0_clk _0021_ VGND VGND VPWR VPWR ram\[29\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold92 ram\[21\]\[6\] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 ram\[36\]\[4\] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 ram\[37\]\[2\] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_18_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2830_ _1085_ net445 _1377_ VGND VGND VPWR VPWR _1384_ sky130_fd_sc_hd__mux2_1
X_2761_ _1087_ net280 _1338_ VGND VGND VPWR VPWR _1346_ sky130_fd_sc_hd__mux2_1
X_2692_ net91 _1188_ _1303_ VGND VGND VPWR VPWR _1306_ sky130_fd_sc_hd__mux2_1
XANTENNA_1 _1048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3313_ _1548_ net234 _1646_ VGND VGND VPWR VPWR _1652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3244_ _1615_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_69_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3175_ _1548_ net431 _1572_ VGND VGND VPWR VPWR _1578_ sky130_fd_sc_hd__mux2_1
X_2126_ ram\[6\]\[5\] ram\[7\]\[5\] _0608_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2057_ ram\[4\]\[4\] ram\[5\]\[4\] _0615_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2959_ _1406_ net200 _1452_ VGND VGND VPWR VPWR _1458_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3931_ clknet_leaf_32_clk _0487_ VGND VGND VPWR VPWR ram\[63\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_3862_ clknet_leaf_34_clk _0424_ VGND VGND VPWR VPWR ram\[57\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2813_ _1374_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3793_ clknet_leaf_25_clk _0355_ VGND VGND VPWR VPWR ram\[48\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2744_ _1087_ net268 _1329_ VGND VGND VPWR VPWR _1337_ sky130_fd_sc_hd__mux2_1
X_2675_ _1077_ net498 _1294_ VGND VGND VPWR VPWR _1297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3227_ _1606_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__clkbuf_1
X_3158_ _1548_ net414 _1563_ VGND VGND VPWR VPWR _1569_ sky130_fd_sc_hd__mux2_1
X_2109_ _0596_ _0903_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__and2_1
X_3089_ _1395_ ram\[50\]\[0\] _1528_ VGND VGND VPWR VPWR _1529_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold381 ram\[29\]\[6\] VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold370 ram\[30\]\[5\] VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 ram\[51\]\[3\] VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2460_ _1176_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__clkbuf_1
X_2391_ _1087_ net206 _1128_ VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_79_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3012_ _1486_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3914_ clknet_leaf_12_clk _0470_ VGND VGND VPWR VPWR ram\[9\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3845_ clknet_leaf_30_clk _0407_ VGND VGND VPWR VPWR ram\[55\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3776_ clknet_leaf_22_clk _0338_ VGND VGND VPWR VPWR ram\[46\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2727_ net378 _1327_ _1313_ VGND VGND VPWR VPWR _1328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2658_ net261 _1188_ _1285_ VGND VGND VPWR VPWR _1288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2589_ _1077_ net123 _1248_ VGND VGND VPWR VPWR _1251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1960_ _0604_ ram\[8\]\[2\] VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__and2b_1
X_1891_ _0614_ _0689_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3630_ clknet_leaf_7_clk _0192_ VGND VGND VPWR VPWR ram\[28\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3561_ clknet_leaf_37_clk _0123_ VGND VGND VPWR VPWR ram\[1\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2512_ _1209_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3492_ clknet_leaf_10_clk _0054_ VGND VGND VPWR VPWR ram\[11\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2443_ _1081_ net230 _1162_ VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__mux2_1
X_2374_ _0535_ _0533_ net15 _0530_ VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_39_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3828_ clknet_leaf_31_clk _0390_ VGND VGND VPWR VPWR ram\[53\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3759_ clknet_leaf_21_clk _0321_ VGND VGND VPWR VPWR ram\[44\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2090_ _0602_ ram\[37\]\[5\] _0570_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2992_ _1404_ net519 _1471_ VGND VGND VPWR VPWR _1476_ sky130_fd_sc_hd__mux2_1
X_1943_ ram\[56\]\[2\] ram\[57\]\[2\] ram\[58\]\[2\] ram\[59\]\[2\] _0615_ _0553_
+ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3613_ clknet_leaf_0_clk _0175_ VGND VGND VPWR VPWR ram\[26\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1874_ _0543_ _0665_ _0672_ _0581_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__a211o_1
XFILLER_0_3_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3544_ clknet_leaf_38_clk _0106_ VGND VGND VPWR VPWR ram\[17\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3475_ clknet_leaf_39_clk _0037_ VGND VGND VPWR VPWR ram\[0\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2426_ _1156_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2357_ _1116_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__clkbuf_1
X_2288_ _0533_ _0535_ net1 VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__and3b_1
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3260_ net283 net11 _1619_ VGND VGND VPWR VPWR _1624_ sky130_fd_sc_hd__mux2_1
X_3191_ _1586_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__clkbuf_1
X_2211_ _0611_ _0996_ _1003_ _0583_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__a211o_1
XFILLER_0_56_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2142_ _0934_ _0935_ _0621_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2073_ _0866_ _0867_ _0868_ _0618_ _0563_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__o221a_1
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2975_ _1466_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__clkbuf_1
X_1926_ ram\[32\]\[2\] ram\[33\]\[2\] ram\[34\]\[2\] ram\[35\]\[2\] _0576_ _0577_
+ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1857_ _0637_ _0648_ _0656_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1788_ _0567_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__clkbuf_4
X_3527_ clknet_leaf_8_clk _0089_ VGND VGND VPWR VPWR ram\[15\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3458_ clknet_leaf_8_clk _0020_ VGND VGND VPWR VPWR ram\[29\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3389_ _1692_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__clkbuf_1
X_2409_ _1146_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_24_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_33_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_42_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold82 ram\[48\]\[1\] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 ram\[10\]\[5\] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 ram\[41\]\[4\] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 ram\[33\]\[1\] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_18_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_51_Left_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2760_ _1345_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__clkbuf_1
X_2691_ _1305_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_2 _1056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3312_ _1651_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_60_Left_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3243_ _1546_ net131 _1610_ VGND VGND VPWR VPWR _1615_ sky130_fd_sc_hd__mux2_1
X_3174_ _1577_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__clkbuf_1
X_2125_ _0614_ _0919_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__or2_1
X_2056_ _0584_ _0844_ _0851_ _0005_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_52_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2958_ _1457_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__clkbuf_1
X_1909_ _0649_ ram\[24\]\[1\] VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__and2b_1
X_2889_ _1408_ net45 _1412_ VGND VGND VPWR VPWR _1419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3930_ clknet_leaf_33_clk _0486_ VGND VGND VPWR VPWR ram\[63\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3861_ clknet_leaf_34_clk _0423_ VGND VGND VPWR VPWR ram\[57\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3792_ clknet_leaf_25_clk _0354_ VGND VGND VPWR VPWR ram\[48\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2812_ net81 _1325_ _1367_ VGND VGND VPWR VPWR _1374_ sky130_fd_sc_hd__mux2_1
X_2743_ _1336_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2674_ _1296_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3226_ _1546_ net228 _1601_ VGND VGND VPWR VPWR _1606_ sky130_fd_sc_hd__mux2_1
X_3157_ _1568_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__clkbuf_1
X_2108_ ram\[56\]\[5\] ram\[57\]\[5\] ram\[58\]\[5\] ram\[59\]\[5\] _0615_ _0652_
+ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_65_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3088_ _1451_ _1509_ VGND VGND VPWR VPWR _1528_ sky130_fd_sc_hd__nand2_4
XFILLER_0_49_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2039_ _0575_ _0834_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold371 ram\[17\]\[3\] VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold360 ram\[46\]\[1\] VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 ram\[49\]\[4\] VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 ram\[55\]\[0\] VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2390_ _1135_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_79_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3011_ _1406_ net63 _1480_ VGND VGND VPWR VPWR _1486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3913_ clknet_leaf_10_clk _0469_ VGND VGND VPWR VPWR ram\[9\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3844_ clknet_leaf_31_clk _0406_ VGND VGND VPWR VPWR ram\[55\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_34_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3775_ clknet_leaf_21_clk _0337_ VGND VGND VPWR VPWR ram\[46\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2726_ net14 VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__clkbuf_4
X_2657_ _1287_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2588_ _1250_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3209_ net73 _1321_ _1592_ VGND VGND VPWR VPWR _1597_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold190 ram\[36\]\[7\] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1890_ ram\[4\]\[1\] ram\[5\]\[1\] _0615_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3560_ clknet_leaf_39_clk _0122_ VGND VGND VPWR VPWR ram\[1\]\[6\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2511_ net72 _1196_ _1202_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__mux2_1
X_3491_ clknet_leaf_10_clk _0053_ VGND VGND VPWR VPWR ram\[11\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2442_ _1166_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__clkbuf_1
X_2373_ _0540_ _0537_ _1124_ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__and3b_2
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3827_ clknet_leaf_29_clk _0389_ VGND VGND VPWR VPWR ram\[53\]\[1\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3758_ clknet_leaf_20_clk _0320_ VGND VGND VPWR VPWR ram\[44\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2709_ net120 _1315_ _1313_ VGND VGND VPWR VPWR _1316_ sky130_fd_sc_hd__mux2_1
X_3689_ clknet_leaf_13_clk _0251_ VGND VGND VPWR VPWR ram\[35\]\[7\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2991_ _1475_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__clkbuf_1
X_1942_ _0737_ _0738_ _0739_ _0606_ _0585_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1873_ _0669_ _0671_ _0542_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__o21ba_1
X_3612_ clknet_leaf_0_clk _0174_ VGND VGND VPWR VPWR ram\[26\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3543_ clknet_leaf_2_clk _0105_ VGND VGND VPWR VPWR ram\[17\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_3474_ clknet_leaf_42_clk _0036_ VGND VGND VPWR VPWR ram\[0\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2425_ _1083_ net375 _1150_ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2356_ net392 _1048_ _1115_ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__mux2_1
X_2287_ _0540_ net5 _0537_ net15 VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__and4b_2
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2210_ _0998_ _1002_ _0003_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__o21ba_1
X_3190_ _1546_ net69 _1581_ VGND VGND VPWR VPWR _1586_ sky130_fd_sc_hd__mux2_1
X_2141_ ram\[30\]\[6\] ram\[31\]\[6\] _0654_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__mux2_1
X_2072_ ram\[10\]\[4\] ram\[11\]\[4\] _0576_ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2974_ _1404_ net508 _1461_ VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__mux2_1
X_1925_ _0720_ _0721_ _0722_ _0606_ _0573_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__o221a_1
X_1856_ _0650_ _0653_ _0655_ _0644_ _0645_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1787_ _0585_ _0586_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3526_ clknet_leaf_8_clk _0088_ VGND VGND VPWR VPWR ram\[15\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3457_ clknet_leaf_37_clk _0019_ VGND VGND VPWR VPWR ram\[7\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3388_ _1048_ net447 _1691_ VGND VGND VPWR VPWR _1692_ sky130_fd_sc_hd__mux2_1
X_2408_ net224 _1066_ _1139_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__mux2_1
X_2339_ net177 _1056_ _1104_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold50 ram\[56\]\[4\] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold61 ram\[20\]\[4\] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 ram\[21\]\[3\] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 ram\[37\]\[3\] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 ram\[2\]\[2\] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_18_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2690_ net256 _1186_ _1303_ VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__mux2_1
XANTENNA_3 _1060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3311_ _1546_ net235 _1646_ VGND VGND VPWR VPWR _1651_ sky130_fd_sc_hd__mux2_1
X_3242_ _1614_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__clkbuf_1
X_3173_ _1546_ net229 _1572_ VGND VGND VPWR VPWR _1577_ sky130_fd_sc_hd__mux2_1
X_2124_ ram\[4\]\[5\] ram\[5\]\[5\] _0615_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__mux2_1
X_2055_ _0848_ _0850_ _0542_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_52_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2957_ _1404_ net469 _1452_ VGND VGND VPWR VPWR _1457_ sky130_fd_sc_hd__mux2_1
X_1908_ ram\[28\]\[1\] ram\[29\]\[1\] ram\[30\]\[1\] ram\[31\]\[1\] _0638_ _0628_
+ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__mux4_1
X_2888_ _1418_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1839_ ram\[12\]\[0\] ram\[13\]\[0\] ram\[14\]\[0\] ram\[15\]\[0\] _0638_ _0624_
+ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__mux4_1
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3509_ clknet_leaf_10_clk _0071_ VGND VGND VPWR VPWR ram\[13\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_68_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_67_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_28_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_2
X_3860_ clknet_leaf_35_clk _0422_ VGND VGND VPWR VPWR ram\[57\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3791_ clknet_leaf_27_clk _0353_ VGND VGND VPWR VPWR ram\[48\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2811_ _1373_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2742_ _1085_ net337 _1329_ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2673_ _1075_ net357 _1294_ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3225_ _1605_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__clkbuf_1
X_3156_ _1546_ net223 _1563_ VGND VGND VPWR VPWR _1568_ sky130_fd_sc_hd__mux2_1
X_2107_ _0899_ _0900_ _0901_ _0606_ _0585_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__o221a_1
X_3087_ _1527_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_65_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_19_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2038_ ram\[32\]\[4\] ram\[33\]\[4\] ram\[34\]\[4\] ram\[35\]\[4\] _0576_ _0553_
+ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_37_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold350 ram\[18\]\[4\] VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 ram\[12\]\[7\] VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 ram\[42\]\[1\] VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 ram\[48\]\[0\] VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 ram\[55\]\[5\] VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3010_ _1485_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3912_ clknet_leaf_4_clk _0468_ VGND VGND VPWR VPWR ram\[9\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_34_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3843_ clknet_leaf_29_clk _0405_ VGND VGND VPWR VPWR ram\[55\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3774_ clknet_leaf_20_clk _0336_ VGND VGND VPWR VPWR ram\[46\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2725_ _1326_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2656_ net140 _1186_ _1285_ VGND VGND VPWR VPWR _1287_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_8_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2587_ _1075_ net259 _1248_ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3208_ _1596_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__clkbuf_1
X_3139_ _1546_ net210 _1554_ VGND VGND VPWR VPWR _1559_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold180 ram\[16\]\[0\] VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 ram\[3\]\[3\] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2510_ _1208_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__clkbuf_1
X_3490_ clknet_leaf_10_clk _0052_ VGND VGND VPWR VPWR ram\[11\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2441_ _1079_ net430 _1162_ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__mux2_1
X_2372_ net5 VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_444 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3826_ clknet_leaf_29_clk _0388_ VGND VGND VPWR VPWR ram\[53\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3757_ clknet_leaf_20_clk _0319_ VGND VGND VPWR VPWR ram\[44\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2708_ net8 VGND VGND VPWR VPWR _1315_ sky130_fd_sc_hd__buf_4
X_3688_ clknet_leaf_13_clk _0250_ VGND VGND VPWR VPWR ram\[35\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2639_ net335 _1186_ _1276_ VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2990_ _1402_ net482 _1471_ VGND VGND VPWR VPWR _1475_ sky130_fd_sc_hd__mux2_1
X_1941_ ram\[62\]\[2\] ram\[63\]\[2\] _0604_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1872_ _0575_ _0670_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__and2_1
X_3611_ clknet_leaf_0_clk _0173_ VGND VGND VPWR VPWR ram\[26\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_3542_ clknet_leaf_43_clk _0104_ VGND VGND VPWR VPWR ram\[17\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3473_ clknet_leaf_13_clk _0035_ VGND VGND VPWR VPWR ram\[8\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2424_ _1155_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__clkbuf_1
X_2355_ _1091_ _1114_ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__nor2_4
X_2286_ net7 VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3809_ clknet_leaf_23_clk _0371_ VGND VGND VPWR VPWR ram\[50\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2140_ _0559_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__clkbuf_4
X_2071_ _0641_ ram\[9\]\[4\] _0550_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2973_ _1465_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1924_ ram\[38\]\[2\] ram\[39\]\[2\] _0649_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1855_ ram\[26\]\[0\] ram\[27\]\[0\] _0654_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__mux2_1
X_1786_ ram\[52\]\[0\] ram\[53\]\[0\] ram\[54\]\[0\] ram\[55\]\[0\] _0547_ _0550_
+ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__mux4_1
X_3525_ clknet_leaf_10_clk _0087_ VGND VGND VPWR VPWR ram\[15\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_3456_ clknet_leaf_37_clk _0018_ VGND VGND VPWR VPWR ram\[7\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3387_ _1441_ _1509_ VGND VGND VPWR VPWR _1691_ sky130_fd_sc_hd__nand2_4
X_2407_ _1145_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__clkbuf_1
X_2338_ _1105_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__clkbuf_1
X_2269_ net363 _1058_ _1054_ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold40 ram\[45\]\[5\] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 ram\[18\]\[6\] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 ram\[4\]\[1\] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 ram\[53\]\[2\] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 ram\[28\]\[0\] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 ram\[9\]\[3\] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_18_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_4 _1081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3310_ _1650_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3241_ _1544_ net168 _1610_ VGND VGND VPWR VPWR _1614_ sky130_fd_sc_hd__mux2_1
X_3172_ _1576_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__clkbuf_1
X_2123_ _0914_ _0916_ _0917_ _0564_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__a22o_1
X_2054_ _0596_ _0849_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2956_ _1456_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__clkbuf_1
X_2887_ _1406_ net369 _1412_ VGND VGND VPWR VPWR _1418_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1907_ _0637_ _0701_ _0705_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1838_ _0567_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__buf_4
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1769_ _0568_ ram\[36\]\[0\] VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__and2b_1
X_3508_ clknet_leaf_9_clk _0070_ VGND VGND VPWR VPWR ram\[13\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3439_ _1718_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_68_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3790_ clknet_leaf_36_clk _0352_ VGND VGND VPWR VPWR ram\[48\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2810_ net56 _1323_ _1367_ VGND VGND VPWR VPWR _1373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2741_ _1335_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2672_ _1295_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3224_ _1544_ net80 _1601_ VGND VGND VPWR VPWR _1605_ sky130_fd_sc_hd__mux2_1
.ends

