magic
tech sky130A
magscale 1 2
timestamp 1703415176
<< obsli1 >>
rect 1104 2159 46092 46801
<< obsm1 >>
rect 1104 2128 46170 46832
<< metal2 >>
rect 22558 48620 22614 49420
rect 25778 48620 25834 49420
rect 27710 48620 27766 49420
rect 28354 48620 28410 49420
rect 14830 0 14886 800
rect 16118 0 16174 800
rect 17406 0 17462 800
rect 19982 0 20038 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
<< obsm2 >>
rect 1400 48564 22502 48620
rect 22670 48564 25722 48620
rect 25890 48564 27654 48620
rect 27822 48564 28298 48620
rect 28466 48564 46166 48620
rect 1400 856 46166 48564
rect 1400 800 14774 856
rect 14942 800 16062 856
rect 16230 800 17350 856
rect 17518 800 19926 856
rect 20094 800 21214 856
rect 21382 800 21858 856
rect 22026 800 22502 856
rect 22670 800 23146 856
rect 23314 800 46166 856
<< metal3 >>
rect 0 45568 800 45688
rect 46476 29248 47276 29368
rect 46476 28568 47276 28688
rect 46476 27888 47276 28008
rect 46476 27208 47276 27328
rect 46476 26528 47276 26648
rect 46476 25848 47276 25968
rect 46476 25168 47276 25288
rect 46476 24488 47276 24608
rect 46476 23808 47276 23928
rect 46476 23128 47276 23248
rect 46476 19048 47276 19168
<< obsm3 >>
rect 800 45768 46476 46817
rect 880 45488 46476 45768
rect 800 29448 46476 45488
rect 800 29168 46396 29448
rect 800 28768 46476 29168
rect 800 28488 46396 28768
rect 800 28088 46476 28488
rect 800 27808 46396 28088
rect 800 27408 46476 27808
rect 800 27128 46396 27408
rect 800 26728 46476 27128
rect 800 26448 46396 26728
rect 800 26048 46476 26448
rect 800 25768 46396 26048
rect 800 25368 46476 25768
rect 800 25088 46396 25368
rect 800 24688 46476 25088
rect 800 24408 46396 24688
rect 800 24008 46476 24408
rect 800 23728 46396 24008
rect 800 23328 46476 23728
rect 800 23048 46396 23328
rect 800 19248 46476 23048
rect 800 18968 46396 19248
rect 800 2143 46476 18968
<< metal4 >>
rect 4208 2128 4528 46832
rect 4868 2128 5188 46832
rect 34928 2128 35248 46832
rect 35588 2128 35908 46832
<< obsm4 >>
rect 11651 2619 34848 42533
rect 35328 2619 35508 42533
rect 35988 2619 40605 42533
<< metal5 >>
rect 1056 36642 46140 36962
rect 1056 35982 46140 36302
rect 1056 6006 46140 6326
rect 1056 5346 46140 5666
<< labels >>
rlabel metal4 s 4868 2128 5188 46832 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 35588 2128 35908 46832 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6006 46140 6326 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 36642 46140 36962 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 46832 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 46832 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5346 46140 5666 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 35982 46140 36302 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 22558 0 22614 800 6 addr[0]
port 3 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 addr[1]
port 4 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 addr[2]
port 5 nsew signal input
rlabel metal2 s 22558 48620 22614 49420 6 addr[3]
port 6 nsew signal input
rlabel metal2 s 25778 48620 25834 49420 6 addr[4]
port 7 nsew signal input
rlabel metal3 s 46476 23808 47276 23928 6 addr[5]
port 8 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 clk
port 9 nsew signal input
rlabel metal2 s 27710 48620 27766 49420 6 data[0]
port 10 nsew signal input
rlabel metal2 s 28354 48620 28410 49420 6 data[1]
port 11 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 data[2]
port 12 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 data[3]
port 13 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 data[4]
port 14 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 data[5]
port 15 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 data[6]
port 16 nsew signal input
rlabel metal3 s 46476 19048 47276 19168 6 data[7]
port 17 nsew signal input
rlabel metal3 s 46476 29248 47276 29368 6 q[0]
port 18 nsew signal output
rlabel metal3 s 46476 25168 47276 25288 6 q[1]
port 19 nsew signal output
rlabel metal3 s 46476 28568 47276 28688 6 q[2]
port 20 nsew signal output
rlabel metal3 s 46476 27888 47276 28008 6 q[3]
port 21 nsew signal output
rlabel metal3 s 46476 27208 47276 27328 6 q[4]
port 22 nsew signal output
rlabel metal3 s 46476 24488 47276 24608 6 q[5]
port 23 nsew signal output
rlabel metal3 s 46476 25848 47276 25968 6 q[6]
port 24 nsew signal output
rlabel metal3 s 46476 26528 47276 26648 6 q[7]
port 25 nsew signal output
rlabel metal3 s 46476 23128 47276 23248 6 we
port 26 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 47276 49420
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6281662
string GDS_FILE /openlane/designs/ram/runs/RUN_2023.12.24_10.45.30/results/signoff/single_port_ram.magic.gds
string GDS_START 393026
<< end >>

