// This is the unpowered netlist.
module single_port_ram (clk,
    we,
    addr,
    data,
    q);
 input clk;
 input we;
 input [5:0] addr;
 input [7:0] data;
 output [7:0] q;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire \addr_reg[0] ;
 wire \addr_reg[1] ;
 wire \addr_reg[2] ;
 wire \addr_reg[3] ;
 wire \addr_reg[4] ;
 wire \addr_reg[5] ;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \ram[0][0] ;
 wire \ram[0][1] ;
 wire \ram[0][2] ;
 wire \ram[0][3] ;
 wire \ram[0][4] ;
 wire \ram[0][5] ;
 wire \ram[0][6] ;
 wire \ram[0][7] ;
 wire \ram[10][0] ;
 wire \ram[10][1] ;
 wire \ram[10][2] ;
 wire \ram[10][3] ;
 wire \ram[10][4] ;
 wire \ram[10][5] ;
 wire \ram[10][6] ;
 wire \ram[10][7] ;
 wire \ram[11][0] ;
 wire \ram[11][1] ;
 wire \ram[11][2] ;
 wire \ram[11][3] ;
 wire \ram[11][4] ;
 wire \ram[11][5] ;
 wire \ram[11][6] ;
 wire \ram[11][7] ;
 wire \ram[12][0] ;
 wire \ram[12][1] ;
 wire \ram[12][2] ;
 wire \ram[12][3] ;
 wire \ram[12][4] ;
 wire \ram[12][5] ;
 wire \ram[12][6] ;
 wire \ram[12][7] ;
 wire \ram[13][0] ;
 wire \ram[13][1] ;
 wire \ram[13][2] ;
 wire \ram[13][3] ;
 wire \ram[13][4] ;
 wire \ram[13][5] ;
 wire \ram[13][6] ;
 wire \ram[13][7] ;
 wire \ram[14][0] ;
 wire \ram[14][1] ;
 wire \ram[14][2] ;
 wire \ram[14][3] ;
 wire \ram[14][4] ;
 wire \ram[14][5] ;
 wire \ram[14][6] ;
 wire \ram[14][7] ;
 wire \ram[15][0] ;
 wire \ram[15][1] ;
 wire \ram[15][2] ;
 wire \ram[15][3] ;
 wire \ram[15][4] ;
 wire \ram[15][5] ;
 wire \ram[15][6] ;
 wire \ram[15][7] ;
 wire \ram[16][0] ;
 wire \ram[16][1] ;
 wire \ram[16][2] ;
 wire \ram[16][3] ;
 wire \ram[16][4] ;
 wire \ram[16][5] ;
 wire \ram[16][6] ;
 wire \ram[16][7] ;
 wire \ram[17][0] ;
 wire \ram[17][1] ;
 wire \ram[17][2] ;
 wire \ram[17][3] ;
 wire \ram[17][4] ;
 wire \ram[17][5] ;
 wire \ram[17][6] ;
 wire \ram[17][7] ;
 wire \ram[18][0] ;
 wire \ram[18][1] ;
 wire \ram[18][2] ;
 wire \ram[18][3] ;
 wire \ram[18][4] ;
 wire \ram[18][5] ;
 wire \ram[18][6] ;
 wire \ram[18][7] ;
 wire \ram[19][0] ;
 wire \ram[19][1] ;
 wire \ram[19][2] ;
 wire \ram[19][3] ;
 wire \ram[19][4] ;
 wire \ram[19][5] ;
 wire \ram[19][6] ;
 wire \ram[19][7] ;
 wire \ram[1][0] ;
 wire \ram[1][1] ;
 wire \ram[1][2] ;
 wire \ram[1][3] ;
 wire \ram[1][4] ;
 wire \ram[1][5] ;
 wire \ram[1][6] ;
 wire \ram[1][7] ;
 wire \ram[20][0] ;
 wire \ram[20][1] ;
 wire \ram[20][2] ;
 wire \ram[20][3] ;
 wire \ram[20][4] ;
 wire \ram[20][5] ;
 wire \ram[20][6] ;
 wire \ram[20][7] ;
 wire \ram[21][0] ;
 wire \ram[21][1] ;
 wire \ram[21][2] ;
 wire \ram[21][3] ;
 wire \ram[21][4] ;
 wire \ram[21][5] ;
 wire \ram[21][6] ;
 wire \ram[21][7] ;
 wire \ram[22][0] ;
 wire \ram[22][1] ;
 wire \ram[22][2] ;
 wire \ram[22][3] ;
 wire \ram[22][4] ;
 wire \ram[22][5] ;
 wire \ram[22][6] ;
 wire \ram[22][7] ;
 wire \ram[23][0] ;
 wire \ram[23][1] ;
 wire \ram[23][2] ;
 wire \ram[23][3] ;
 wire \ram[23][4] ;
 wire \ram[23][5] ;
 wire \ram[23][6] ;
 wire \ram[23][7] ;
 wire \ram[24][0] ;
 wire \ram[24][1] ;
 wire \ram[24][2] ;
 wire \ram[24][3] ;
 wire \ram[24][4] ;
 wire \ram[24][5] ;
 wire \ram[24][6] ;
 wire \ram[24][7] ;
 wire \ram[25][0] ;
 wire \ram[25][1] ;
 wire \ram[25][2] ;
 wire \ram[25][3] ;
 wire \ram[25][4] ;
 wire \ram[25][5] ;
 wire \ram[25][6] ;
 wire \ram[25][7] ;
 wire \ram[26][0] ;
 wire \ram[26][1] ;
 wire \ram[26][2] ;
 wire \ram[26][3] ;
 wire \ram[26][4] ;
 wire \ram[26][5] ;
 wire \ram[26][6] ;
 wire \ram[26][7] ;
 wire \ram[27][0] ;
 wire \ram[27][1] ;
 wire \ram[27][2] ;
 wire \ram[27][3] ;
 wire \ram[27][4] ;
 wire \ram[27][5] ;
 wire \ram[27][6] ;
 wire \ram[27][7] ;
 wire \ram[28][0] ;
 wire \ram[28][1] ;
 wire \ram[28][2] ;
 wire \ram[28][3] ;
 wire \ram[28][4] ;
 wire \ram[28][5] ;
 wire \ram[28][6] ;
 wire \ram[28][7] ;
 wire \ram[29][0] ;
 wire \ram[29][1] ;
 wire \ram[29][2] ;
 wire \ram[29][3] ;
 wire \ram[29][4] ;
 wire \ram[29][5] ;
 wire \ram[29][6] ;
 wire \ram[29][7] ;
 wire \ram[2][0] ;
 wire \ram[2][1] ;
 wire \ram[2][2] ;
 wire \ram[2][3] ;
 wire \ram[2][4] ;
 wire \ram[2][5] ;
 wire \ram[2][6] ;
 wire \ram[2][7] ;
 wire \ram[30][0] ;
 wire \ram[30][1] ;
 wire \ram[30][2] ;
 wire \ram[30][3] ;
 wire \ram[30][4] ;
 wire \ram[30][5] ;
 wire \ram[30][6] ;
 wire \ram[30][7] ;
 wire \ram[31][0] ;
 wire \ram[31][1] ;
 wire \ram[31][2] ;
 wire \ram[31][3] ;
 wire \ram[31][4] ;
 wire \ram[31][5] ;
 wire \ram[31][6] ;
 wire \ram[31][7] ;
 wire \ram[32][0] ;
 wire \ram[32][1] ;
 wire \ram[32][2] ;
 wire \ram[32][3] ;
 wire \ram[32][4] ;
 wire \ram[32][5] ;
 wire \ram[32][6] ;
 wire \ram[32][7] ;
 wire \ram[33][0] ;
 wire \ram[33][1] ;
 wire \ram[33][2] ;
 wire \ram[33][3] ;
 wire \ram[33][4] ;
 wire \ram[33][5] ;
 wire \ram[33][6] ;
 wire \ram[33][7] ;
 wire \ram[34][0] ;
 wire \ram[34][1] ;
 wire \ram[34][2] ;
 wire \ram[34][3] ;
 wire \ram[34][4] ;
 wire \ram[34][5] ;
 wire \ram[34][6] ;
 wire \ram[34][7] ;
 wire \ram[35][0] ;
 wire \ram[35][1] ;
 wire \ram[35][2] ;
 wire \ram[35][3] ;
 wire \ram[35][4] ;
 wire \ram[35][5] ;
 wire \ram[35][6] ;
 wire \ram[35][7] ;
 wire \ram[36][0] ;
 wire \ram[36][1] ;
 wire \ram[36][2] ;
 wire \ram[36][3] ;
 wire \ram[36][4] ;
 wire \ram[36][5] ;
 wire \ram[36][6] ;
 wire \ram[36][7] ;
 wire \ram[37][0] ;
 wire \ram[37][1] ;
 wire \ram[37][2] ;
 wire \ram[37][3] ;
 wire \ram[37][4] ;
 wire \ram[37][5] ;
 wire \ram[37][6] ;
 wire \ram[37][7] ;
 wire \ram[38][0] ;
 wire \ram[38][1] ;
 wire \ram[38][2] ;
 wire \ram[38][3] ;
 wire \ram[38][4] ;
 wire \ram[38][5] ;
 wire \ram[38][6] ;
 wire \ram[38][7] ;
 wire \ram[39][0] ;
 wire \ram[39][1] ;
 wire \ram[39][2] ;
 wire \ram[39][3] ;
 wire \ram[39][4] ;
 wire \ram[39][5] ;
 wire \ram[39][6] ;
 wire \ram[39][7] ;
 wire \ram[3][0] ;
 wire \ram[3][1] ;
 wire \ram[3][2] ;
 wire \ram[3][3] ;
 wire \ram[3][4] ;
 wire \ram[3][5] ;
 wire \ram[3][6] ;
 wire \ram[3][7] ;
 wire \ram[40][0] ;
 wire \ram[40][1] ;
 wire \ram[40][2] ;
 wire \ram[40][3] ;
 wire \ram[40][4] ;
 wire \ram[40][5] ;
 wire \ram[40][6] ;
 wire \ram[40][7] ;
 wire \ram[41][0] ;
 wire \ram[41][1] ;
 wire \ram[41][2] ;
 wire \ram[41][3] ;
 wire \ram[41][4] ;
 wire \ram[41][5] ;
 wire \ram[41][6] ;
 wire \ram[41][7] ;
 wire \ram[42][0] ;
 wire \ram[42][1] ;
 wire \ram[42][2] ;
 wire \ram[42][3] ;
 wire \ram[42][4] ;
 wire \ram[42][5] ;
 wire \ram[42][6] ;
 wire \ram[42][7] ;
 wire \ram[43][0] ;
 wire \ram[43][1] ;
 wire \ram[43][2] ;
 wire \ram[43][3] ;
 wire \ram[43][4] ;
 wire \ram[43][5] ;
 wire \ram[43][6] ;
 wire \ram[43][7] ;
 wire \ram[44][0] ;
 wire \ram[44][1] ;
 wire \ram[44][2] ;
 wire \ram[44][3] ;
 wire \ram[44][4] ;
 wire \ram[44][5] ;
 wire \ram[44][6] ;
 wire \ram[44][7] ;
 wire \ram[45][0] ;
 wire \ram[45][1] ;
 wire \ram[45][2] ;
 wire \ram[45][3] ;
 wire \ram[45][4] ;
 wire \ram[45][5] ;
 wire \ram[45][6] ;
 wire \ram[45][7] ;
 wire \ram[46][0] ;
 wire \ram[46][1] ;
 wire \ram[46][2] ;
 wire \ram[46][3] ;
 wire \ram[46][4] ;
 wire \ram[46][5] ;
 wire \ram[46][6] ;
 wire \ram[46][7] ;
 wire \ram[47][0] ;
 wire \ram[47][1] ;
 wire \ram[47][2] ;
 wire \ram[47][3] ;
 wire \ram[47][4] ;
 wire \ram[47][5] ;
 wire \ram[47][6] ;
 wire \ram[47][7] ;
 wire \ram[48][0] ;
 wire \ram[48][1] ;
 wire \ram[48][2] ;
 wire \ram[48][3] ;
 wire \ram[48][4] ;
 wire \ram[48][5] ;
 wire \ram[48][6] ;
 wire \ram[48][7] ;
 wire \ram[49][0] ;
 wire \ram[49][1] ;
 wire \ram[49][2] ;
 wire \ram[49][3] ;
 wire \ram[49][4] ;
 wire \ram[49][5] ;
 wire \ram[49][6] ;
 wire \ram[49][7] ;
 wire \ram[4][0] ;
 wire \ram[4][1] ;
 wire \ram[4][2] ;
 wire \ram[4][3] ;
 wire \ram[4][4] ;
 wire \ram[4][5] ;
 wire \ram[4][6] ;
 wire \ram[4][7] ;
 wire \ram[50][0] ;
 wire \ram[50][1] ;
 wire \ram[50][2] ;
 wire \ram[50][3] ;
 wire \ram[50][4] ;
 wire \ram[50][5] ;
 wire \ram[50][6] ;
 wire \ram[50][7] ;
 wire \ram[51][0] ;
 wire \ram[51][1] ;
 wire \ram[51][2] ;
 wire \ram[51][3] ;
 wire \ram[51][4] ;
 wire \ram[51][5] ;
 wire \ram[51][6] ;
 wire \ram[51][7] ;
 wire \ram[52][0] ;
 wire \ram[52][1] ;
 wire \ram[52][2] ;
 wire \ram[52][3] ;
 wire \ram[52][4] ;
 wire \ram[52][5] ;
 wire \ram[52][6] ;
 wire \ram[52][7] ;
 wire \ram[53][0] ;
 wire \ram[53][1] ;
 wire \ram[53][2] ;
 wire \ram[53][3] ;
 wire \ram[53][4] ;
 wire \ram[53][5] ;
 wire \ram[53][6] ;
 wire \ram[53][7] ;
 wire \ram[54][0] ;
 wire \ram[54][1] ;
 wire \ram[54][2] ;
 wire \ram[54][3] ;
 wire \ram[54][4] ;
 wire \ram[54][5] ;
 wire \ram[54][6] ;
 wire \ram[54][7] ;
 wire \ram[55][0] ;
 wire \ram[55][1] ;
 wire \ram[55][2] ;
 wire \ram[55][3] ;
 wire \ram[55][4] ;
 wire \ram[55][5] ;
 wire \ram[55][6] ;
 wire \ram[55][7] ;
 wire \ram[56][0] ;
 wire \ram[56][1] ;
 wire \ram[56][2] ;
 wire \ram[56][3] ;
 wire \ram[56][4] ;
 wire \ram[56][5] ;
 wire \ram[56][6] ;
 wire \ram[56][7] ;
 wire \ram[57][0] ;
 wire \ram[57][1] ;
 wire \ram[57][2] ;
 wire \ram[57][3] ;
 wire \ram[57][4] ;
 wire \ram[57][5] ;
 wire \ram[57][6] ;
 wire \ram[57][7] ;
 wire \ram[58][0] ;
 wire \ram[58][1] ;
 wire \ram[58][2] ;
 wire \ram[58][3] ;
 wire \ram[58][4] ;
 wire \ram[58][5] ;
 wire \ram[58][6] ;
 wire \ram[58][7] ;
 wire \ram[59][0] ;
 wire \ram[59][1] ;
 wire \ram[59][2] ;
 wire \ram[59][3] ;
 wire \ram[59][4] ;
 wire \ram[59][5] ;
 wire \ram[59][6] ;
 wire \ram[59][7] ;
 wire \ram[5][0] ;
 wire \ram[5][1] ;
 wire \ram[5][2] ;
 wire \ram[5][3] ;
 wire \ram[5][4] ;
 wire \ram[5][5] ;
 wire \ram[5][6] ;
 wire \ram[5][7] ;
 wire \ram[60][0] ;
 wire \ram[60][1] ;
 wire \ram[60][2] ;
 wire \ram[60][3] ;
 wire \ram[60][4] ;
 wire \ram[60][5] ;
 wire \ram[60][6] ;
 wire \ram[60][7] ;
 wire \ram[61][0] ;
 wire \ram[61][1] ;
 wire \ram[61][2] ;
 wire \ram[61][3] ;
 wire \ram[61][4] ;
 wire \ram[61][5] ;
 wire \ram[61][6] ;
 wire \ram[61][7] ;
 wire \ram[62][0] ;
 wire \ram[62][1] ;
 wire \ram[62][2] ;
 wire \ram[62][3] ;
 wire \ram[62][4] ;
 wire \ram[62][5] ;
 wire \ram[62][6] ;
 wire \ram[62][7] ;
 wire \ram[63][0] ;
 wire \ram[63][1] ;
 wire \ram[63][2] ;
 wire \ram[63][3] ;
 wire \ram[63][4] ;
 wire \ram[63][5] ;
 wire \ram[63][6] ;
 wire \ram[63][7] ;
 wire \ram[6][0] ;
 wire \ram[6][1] ;
 wire \ram[6][2] ;
 wire \ram[6][3] ;
 wire \ram[6][4] ;
 wire \ram[6][5] ;
 wire \ram[6][6] ;
 wire \ram[6][7] ;
 wire \ram[7][0] ;
 wire \ram[7][1] ;
 wire \ram[7][2] ;
 wire \ram[7][3] ;
 wire \ram[7][4] ;
 wire \ram[7][5] ;
 wire \ram[7][6] ;
 wire \ram[7][7] ;
 wire \ram[8][0] ;
 wire \ram[8][1] ;
 wire \ram[8][2] ;
 wire \ram[8][3] ;
 wire \ram[8][4] ;
 wire \ram[8][5] ;
 wire \ram[8][6] ;
 wire \ram[8][7] ;
 wire \ram[9][0] ;
 wire \ram[9][1] ;
 wire \ram[9][2] ;
 wire \ram[9][3] ;
 wire \ram[9][4] ;
 wire \ram[9][5] ;
 wire \ram[9][6] ;
 wire \ram[9][7] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_1048_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_1064_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_1056_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_1323_));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_256 ();
 sky130_fd_sc_hd__clkbuf_2 _1724_ (.A(net1),
    .X(_0530_));
 sky130_fd_sc_hd__clkbuf_4 _1725_ (.A(net15),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _1726_ (.A0(_0530_),
    .A1(net463),
    .S(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__clkbuf_1 _1727_ (.A(_0532_),
    .X(_0006_));
 sky130_fd_sc_hd__buf_2 _1728_ (.A(net2),
    .X(_0533_));
 sky130_fd_sc_hd__mux2_1 _1729_ (.A0(_0533_),
    .A1(\addr_reg[1] ),
    .S(_0531_),
    .X(_0534_));
 sky130_fd_sc_hd__clkbuf_1 _1730_ (.A(_0534_),
    .X(_0007_));
 sky130_fd_sc_hd__clkbuf_2 _1731_ (.A(net3),
    .X(_0535_));
 sky130_fd_sc_hd__mux2_1 _1732_ (.A0(_0535_),
    .A1(\addr_reg[2] ),
    .S(_0531_),
    .X(_0536_));
 sky130_fd_sc_hd__clkbuf_1 _1733_ (.A(_0536_),
    .X(_0008_));
 sky130_fd_sc_hd__buf_2 _1734_ (.A(net4),
    .X(_0537_));
 sky130_fd_sc_hd__mux2_1 _1735_ (.A0(_0537_),
    .A1(net197),
    .S(_0531_),
    .X(_0538_));
 sky130_fd_sc_hd__clkbuf_1 _1736_ (.A(_0538_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _1737_ (.A0(net5),
    .A1(net282),
    .S(_0531_),
    .X(_0539_));
 sky130_fd_sc_hd__clkbuf_1 _1738_ (.A(_0539_),
    .X(_0010_));
 sky130_fd_sc_hd__buf_2 _1739_ (.A(net6),
    .X(_0540_));
 sky130_fd_sc_hd__mux2_1 _1740_ (.A0(_0540_),
    .A1(net24),
    .S(_0531_),
    .X(_0541_));
 sky130_fd_sc_hd__clkbuf_1 _1741_ (.A(_0541_),
    .X(_0011_));
 sky130_fd_sc_hd__clkbuf_4 _1742_ (.A(_0003_),
    .X(_0542_));
 sky130_fd_sc_hd__clkbuf_4 _1743_ (.A(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__clkbuf_4 _1744_ (.A(_0002_),
    .X(_0544_));
 sky130_fd_sc_hd__clkbuf_4 _1745_ (.A(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__clkbuf_4 _1746_ (.A(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__buf_4 _1747_ (.A(_0000_),
    .X(_0547_));
 sky130_fd_sc_hd__buf_4 _1748_ (.A(_0547_),
    .X(_0548_));
 sky130_fd_sc_hd__clkbuf_4 _1749_ (.A(_0001_),
    .X(_0549_));
 sky130_fd_sc_hd__buf_4 _1750_ (.A(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__buf_4 _1751_ (.A(_0550_),
    .X(_0551_));
 sky130_fd_sc_hd__mux4_1 _1752_ (.A0(\ram[44][0] ),
    .A1(\ram[45][0] ),
    .A2(\ram[46][0] ),
    .A3(\ram[47][0] ),
    .S0(_0548_),
    .S1(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__buf_4 _1753_ (.A(_0549_),
    .X(_0553_));
 sky130_fd_sc_hd__buf_2 _1754_ (.A(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__clkbuf_4 _1755_ (.A(_0000_),
    .X(_0555_));
 sky130_fd_sc_hd__buf_4 _1756_ (.A(_0555_),
    .X(_0556_));
 sky130_fd_sc_hd__mux2_1 _1757_ (.A0(\ram[40][0] ),
    .A1(\ram[41][0] ),
    .S(_0556_),
    .X(_0557_));
 sky130_fd_sc_hd__or2_1 _1758_ (.A(_0554_),
    .B(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__inv_2 _1759_ (.A(_0001_),
    .Y(_0559_));
 sky130_fd_sc_hd__clkbuf_4 _1760_ (.A(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__clkbuf_8 _1761_ (.A(_0555_),
    .X(_0561_));
 sky130_fd_sc_hd__mux2_1 _1762_ (.A0(\ram[42][0] ),
    .A1(\ram[43][0] ),
    .S(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__clkinv_4 _1763_ (.A(_0002_),
    .Y(_0563_));
 sky130_fd_sc_hd__clkbuf_4 _1764_ (.A(_0563_),
    .X(_0564_));
 sky130_fd_sc_hd__o21a_1 _1765_ (.A1(_0560_),
    .A2(_0562_),
    .B1(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__a22o_1 _1766_ (.A1(_0546_),
    .A2(_0552_),
    .B1(_0558_),
    .B2(_0565_),
    .X(_0566_));
 sky130_fd_sc_hd__buf_4 _1767_ (.A(_0000_),
    .X(_0567_));
 sky130_fd_sc_hd__clkbuf_4 _1768_ (.A(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__and2b_1 _1769_ (.A_N(_0568_),
    .B(\ram[36][0] ),
    .X(_0569_));
 sky130_fd_sc_hd__clkbuf_4 _1770_ (.A(_0549_),
    .X(_0570_));
 sky130_fd_sc_hd__a21o_1 _1771_ (.A1(_0548_),
    .A2(\ram[37][0] ),
    .B1(_0570_),
    .X(_0571_));
 sky130_fd_sc_hd__mux2_1 _1772_ (.A0(\ram[38][0] ),
    .A1(\ram[39][0] ),
    .S(_0556_),
    .X(_0572_));
 sky130_fd_sc_hd__buf_4 _1773_ (.A(_0544_),
    .X(_0573_));
 sky130_fd_sc_hd__o221a_1 _1774_ (.A1(_0569_),
    .A2(_0571_),
    .B1(_0572_),
    .B2(_0560_),
    .C1(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__clkbuf_4 _1775_ (.A(_0563_),
    .X(_0575_));
 sky130_fd_sc_hd__buf_4 _1776_ (.A(_0000_),
    .X(_0576_));
 sky130_fd_sc_hd__buf_4 _1777_ (.A(_0549_),
    .X(_0577_));
 sky130_fd_sc_hd__mux4_1 _1778_ (.A0(\ram[32][0] ),
    .A1(\ram[33][0] ),
    .A2(\ram[34][0] ),
    .A3(\ram[35][0] ),
    .S0(_0576_),
    .S1(_0577_),
    .X(_0578_));
 sky130_fd_sc_hd__and2_1 _1779_ (.A(_0575_),
    .B(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__o21ba_1 _1780_ (.A1(_0574_),
    .A2(_0579_),
    .B1_N(_0542_),
    .X(_0580_));
 sky130_fd_sc_hd__clkbuf_4 _1781_ (.A(_0004_),
    .X(_0581_));
 sky130_fd_sc_hd__a211o_1 _1782_ (.A1(_0543_),
    .A2(_0566_),
    .B1(_0580_),
    .C1(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__inv_2 _1783_ (.A(_0004_),
    .Y(_0583_));
 sky130_fd_sc_hd__clkbuf_4 _1784_ (.A(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__clkbuf_4 _1785_ (.A(_0544_),
    .X(_0585_));
 sky130_fd_sc_hd__mux4_1 _1786_ (.A0(\ram[52][0] ),
    .A1(\ram[53][0] ),
    .A2(\ram[54][0] ),
    .A3(\ram[55][0] ),
    .S0(_0547_),
    .S1(_0550_),
    .X(_0586_));
 sky130_fd_sc_hd__and2_1 _1787_ (.A(_0585_),
    .B(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__clkbuf_4 _1788_ (.A(_0567_),
    .X(_0588_));
 sky130_fd_sc_hd__and2b_1 _1789_ (.A_N(_0588_),
    .B(\ram[48][0] ),
    .X(_0589_));
 sky130_fd_sc_hd__buf_4 _1790_ (.A(_0567_),
    .X(_0590_));
 sky130_fd_sc_hd__clkbuf_4 _1791_ (.A(_0549_),
    .X(_0591_));
 sky130_fd_sc_hd__a21o_1 _1792_ (.A1(_0590_),
    .A2(\ram[49][0] ),
    .B1(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__buf_4 _1793_ (.A(_0555_),
    .X(_0593_));
 sky130_fd_sc_hd__mux2_1 _1794_ (.A0(\ram[50][0] ),
    .A1(\ram[51][0] ),
    .S(_0593_),
    .X(_0594_));
 sky130_fd_sc_hd__clkbuf_4 _1795_ (.A(_0559_),
    .X(_0595_));
 sky130_fd_sc_hd__buf_2 _1796_ (.A(_0563_),
    .X(_0596_));
 sky130_fd_sc_hd__o221a_1 _1797_ (.A1(_0589_),
    .A2(_0592_),
    .B1(_0594_),
    .B2(_0595_),
    .C1(_0596_),
    .X(_0597_));
 sky130_fd_sc_hd__buf_2 _1798_ (.A(_0003_),
    .X(_0598_));
 sky130_fd_sc_hd__o21ba_1 _1799_ (.A1(_0587_),
    .A2(_0597_),
    .B1_N(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__buf_4 _1800_ (.A(_0567_),
    .X(_0600_));
 sky130_fd_sc_hd__and2b_1 _1801_ (.A_N(_0600_),
    .B(\ram[60][0] ),
    .X(_0601_));
 sky130_fd_sc_hd__buf_4 _1802_ (.A(_0547_),
    .X(_0602_));
 sky130_fd_sc_hd__a21o_1 _1803_ (.A1(_0602_),
    .A2(\ram[61][0] ),
    .B1(_0570_),
    .X(_0603_));
 sky130_fd_sc_hd__buf_4 _1804_ (.A(_0555_),
    .X(_0604_));
 sky130_fd_sc_hd__mux2_1 _1805_ (.A0(\ram[62][0] ),
    .A1(\ram[63][0] ),
    .S(_0604_),
    .X(_0605_));
 sky130_fd_sc_hd__clkbuf_4 _1806_ (.A(_0559_),
    .X(_0606_));
 sky130_fd_sc_hd__o221a_1 _1807_ (.A1(_0601_),
    .A2(_0603_),
    .B1(_0605_),
    .B2(_0606_),
    .C1(_0573_),
    .X(_0607_));
 sky130_fd_sc_hd__clkbuf_8 _1808_ (.A(_0000_),
    .X(_0608_));
 sky130_fd_sc_hd__mux4_1 _1809_ (.A0(\ram[56][0] ),
    .A1(\ram[57][0] ),
    .A2(\ram[58][0] ),
    .A3(\ram[59][0] ),
    .S0(_0608_),
    .S1(_0553_),
    .X(_0609_));
 sky130_fd_sc_hd__and2_1 _1810_ (.A(_0575_),
    .B(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__buf_4 _1811_ (.A(_0003_),
    .X(_0611_));
 sky130_fd_sc_hd__o21a_1 _1812_ (.A1(_0607_),
    .A2(_0610_),
    .B1(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__o31a_1 _1813_ (.A1(_0584_),
    .A2(_0599_),
    .A3(_0612_),
    .B1(_0005_),
    .X(_0613_));
 sky130_fd_sc_hd__clkbuf_4 _1814_ (.A(_0549_),
    .X(_0614_));
 sky130_fd_sc_hd__buf_4 _1815_ (.A(_0000_),
    .X(_0615_));
 sky130_fd_sc_hd__mux2_1 _1816_ (.A0(\ram[4][0] ),
    .A1(\ram[5][0] ),
    .S(_0615_),
    .X(_0616_));
 sky130_fd_sc_hd__or2_1 _1817_ (.A(_0614_),
    .B(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__clkbuf_4 _1818_ (.A(_0559_),
    .X(_0618_));
 sky130_fd_sc_hd__buf_4 _1819_ (.A(_0555_),
    .X(_0619_));
 sky130_fd_sc_hd__mux2_1 _1820_ (.A0(\ram[6][0] ),
    .A1(\ram[7][0] ),
    .S(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__clkbuf_4 _1821_ (.A(_0544_),
    .X(_0621_));
 sky130_fd_sc_hd__o21a_1 _1822_ (.A1(_0618_),
    .A2(_0620_),
    .B1(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__buf_4 _1823_ (.A(_0567_),
    .X(_0623_));
 sky130_fd_sc_hd__buf_4 _1824_ (.A(_0549_),
    .X(_0624_));
 sky130_fd_sc_hd__mux4_1 _1825_ (.A0(\ram[0][0] ),
    .A1(\ram[1][0] ),
    .A2(\ram[2][0] ),
    .A3(\ram[3][0] ),
    .S0(_0623_),
    .S1(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__clkbuf_4 _1826_ (.A(_0563_),
    .X(_0626_));
 sky130_fd_sc_hd__a22o_1 _1827_ (.A1(_0617_),
    .A2(_0622_),
    .B1(_0625_),
    .B2(_0626_),
    .X(_0627_));
 sky130_fd_sc_hd__buf_2 _1828_ (.A(_0549_),
    .X(_0628_));
 sky130_fd_sc_hd__buf_4 _1829_ (.A(_0000_),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _1830_ (.A0(\ram[20][0] ),
    .A1(\ram[21][0] ),
    .S(_0629_),
    .X(_0630_));
 sky130_fd_sc_hd__or2_1 _1831_ (.A(_0628_),
    .B(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__mux2_1 _1832_ (.A0(\ram[22][0] ),
    .A1(\ram[23][0] ),
    .S(_0608_),
    .X(_0632_));
 sky130_fd_sc_hd__o21a_1 _1833_ (.A1(_0618_),
    .A2(_0632_),
    .B1(_0544_),
    .X(_0633_));
 sky130_fd_sc_hd__buf_4 _1834_ (.A(_0549_),
    .X(_0634_));
 sky130_fd_sc_hd__mux4_2 _1835_ (.A0(\ram[16][0] ),
    .A1(\ram[17][0] ),
    .A2(\ram[18][0] ),
    .A3(\ram[19][0] ),
    .S0(_0588_),
    .S1(_0634_),
    .X(_0635_));
 sky130_fd_sc_hd__a22o_1 _1836_ (.A1(_0631_),
    .A2(_0633_),
    .B1(_0635_),
    .B2(_0626_),
    .X(_0636_));
 sky130_fd_sc_hd__clkbuf_4 _1837_ (.A(_0545_),
    .X(_0637_));
 sky130_fd_sc_hd__buf_4 _1838_ (.A(_0567_),
    .X(_0638_));
 sky130_fd_sc_hd__mux4_1 _1839_ (.A0(\ram[12][0] ),
    .A1(\ram[13][0] ),
    .A2(\ram[14][0] ),
    .A3(\ram[15][0] ),
    .S0(_0638_),
    .S1(_0624_),
    .X(_0639_));
 sky130_fd_sc_hd__and2b_1 _1840_ (.A_N(_0604_),
    .B(\ram[8][0] ),
    .X(_0640_));
 sky130_fd_sc_hd__clkbuf_4 _1841_ (.A(_0555_),
    .X(_0641_));
 sky130_fd_sc_hd__a21o_1 _1842_ (.A1(_0641_),
    .A2(\ram[9][0] ),
    .B1(_0550_),
    .X(_0642_));
 sky130_fd_sc_hd__mux2_1 _1843_ (.A0(\ram[10][0] ),
    .A1(\ram[11][0] ),
    .S(_0576_),
    .X(_0643_));
 sky130_fd_sc_hd__clkbuf_4 _1844_ (.A(_0559_),
    .X(_0644_));
 sky130_fd_sc_hd__buf_4 _1845_ (.A(_0563_),
    .X(_0645_));
 sky130_fd_sc_hd__o221a_1 _1846_ (.A1(_0640_),
    .A2(_0642_),
    .B1(_0643_),
    .B2(_0644_),
    .C1(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__a21o_1 _1847_ (.A1(_0637_),
    .A2(_0639_),
    .B1(_0646_),
    .X(_0647_));
 sky130_fd_sc_hd__mux4_1 _1848_ (.A0(\ram[28][0] ),
    .A1(\ram[29][0] ),
    .A2(\ram[30][0] ),
    .A3(\ram[31][0] ),
    .S0(_0638_),
    .S1(_0628_),
    .X(_0648_));
 sky130_fd_sc_hd__buf_4 _1849_ (.A(_0555_),
    .X(_0649_));
 sky130_fd_sc_hd__and2b_1 _1850_ (.A_N(_0649_),
    .B(\ram[24][0] ),
    .X(_0650_));
 sky130_fd_sc_hd__buf_4 _1851_ (.A(_0555_),
    .X(_0651_));
 sky130_fd_sc_hd__buf_4 _1852_ (.A(_0549_),
    .X(_0652_));
 sky130_fd_sc_hd__a21o_1 _1853_ (.A1(_0651_),
    .A2(\ram[25][0] ),
    .B1(_0652_),
    .X(_0653_));
 sky130_fd_sc_hd__buf_4 _1854_ (.A(_0555_),
    .X(_0654_));
 sky130_fd_sc_hd__mux2_1 _1855_ (.A0(\ram[26][0] ),
    .A1(\ram[27][0] ),
    .S(_0654_),
    .X(_0655_));
 sky130_fd_sc_hd__o221a_1 _1856_ (.A1(_0650_),
    .A2(_0653_),
    .B1(_0655_),
    .B2(_0644_),
    .C1(_0645_),
    .X(_0656_));
 sky130_fd_sc_hd__a21o_1 _1857_ (.A1(_0637_),
    .A2(_0648_),
    .B1(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__mux4_2 _1858_ (.A0(_0627_),
    .A1(_0636_),
    .A2(_0647_),
    .A3(_0657_),
    .S0(_0004_),
    .S1(_0543_),
    .X(_0658_));
 sky130_fd_sc_hd__inv_2 _1859_ (.A(_0005_),
    .Y(_0659_));
 sky130_fd_sc_hd__a22o_1 _1860_ (.A1(_0582_),
    .A2(_0613_),
    .B1(_0658_),
    .B2(_0659_),
    .X(net16));
 sky130_fd_sc_hd__mux4_1 _1861_ (.A0(\ram[44][1] ),
    .A1(\ram[45][1] ),
    .A2(\ram[46][1] ),
    .A3(\ram[47][1] ),
    .S0(_0548_),
    .S1(_0551_),
    .X(_0660_));
 sky130_fd_sc_hd__mux2_1 _1862_ (.A0(\ram[40][1] ),
    .A1(\ram[41][1] ),
    .S(_0556_),
    .X(_0661_));
 sky130_fd_sc_hd__or2_1 _1863_ (.A(_0554_),
    .B(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__mux2_1 _1864_ (.A0(\ram[42][1] ),
    .A1(\ram[43][1] ),
    .S(_0561_),
    .X(_0663_));
 sky130_fd_sc_hd__o21a_1 _1865_ (.A1(_0560_),
    .A2(_0663_),
    .B1(_0564_),
    .X(_0664_));
 sky130_fd_sc_hd__a22o_1 _1866_ (.A1(_0546_),
    .A2(_0660_),
    .B1(_0662_),
    .B2(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__and2b_1 _1867_ (.A_N(_0568_),
    .B(\ram[36][1] ),
    .X(_0666_));
 sky130_fd_sc_hd__a21o_1 _1868_ (.A1(_0548_),
    .A2(\ram[37][1] ),
    .B1(_0570_),
    .X(_0667_));
 sky130_fd_sc_hd__mux2_1 _1869_ (.A0(\ram[38][1] ),
    .A1(\ram[39][1] ),
    .S(_0556_),
    .X(_0668_));
 sky130_fd_sc_hd__o221a_1 _1870_ (.A1(_0666_),
    .A2(_0667_),
    .B1(_0668_),
    .B2(_0560_),
    .C1(_0573_),
    .X(_0669_));
 sky130_fd_sc_hd__mux4_1 _1871_ (.A0(\ram[32][1] ),
    .A1(\ram[33][1] ),
    .A2(\ram[34][1] ),
    .A3(\ram[35][1] ),
    .S0(_0576_),
    .S1(_0577_),
    .X(_0670_));
 sky130_fd_sc_hd__and2_1 _1872_ (.A(_0575_),
    .B(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__o21ba_1 _1873_ (.A1(_0669_),
    .A2(_0671_),
    .B1_N(_0542_),
    .X(_0672_));
 sky130_fd_sc_hd__a211o_1 _1874_ (.A1(_0543_),
    .A2(_0665_),
    .B1(_0672_),
    .C1(_0581_),
    .X(_0673_));
 sky130_fd_sc_hd__mux4_1 _1875_ (.A0(\ram[52][1] ),
    .A1(\ram[53][1] ),
    .A2(\ram[54][1] ),
    .A3(\ram[55][1] ),
    .S0(_0547_),
    .S1(_0550_),
    .X(_0674_));
 sky130_fd_sc_hd__and2_1 _1876_ (.A(_0585_),
    .B(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__and2b_1 _1877_ (.A_N(_0588_),
    .B(\ram[48][1] ),
    .X(_0676_));
 sky130_fd_sc_hd__a21o_1 _1878_ (.A1(_0590_),
    .A2(\ram[49][1] ),
    .B1(_0591_),
    .X(_0677_));
 sky130_fd_sc_hd__mux2_1 _1879_ (.A0(\ram[50][1] ),
    .A1(\ram[51][1] ),
    .S(_0593_),
    .X(_0678_));
 sky130_fd_sc_hd__o221a_1 _1880_ (.A1(_0676_),
    .A2(_0677_),
    .B1(_0678_),
    .B2(_0595_),
    .C1(_0596_),
    .X(_0679_));
 sky130_fd_sc_hd__o21ba_1 _1881_ (.A1(_0675_),
    .A2(_0679_),
    .B1_N(_0598_),
    .X(_0680_));
 sky130_fd_sc_hd__and2b_1 _1882_ (.A_N(_0600_),
    .B(\ram[60][1] ),
    .X(_0681_));
 sky130_fd_sc_hd__a21o_1 _1883_ (.A1(_0602_),
    .A2(\ram[61][1] ),
    .B1(_0570_),
    .X(_0682_));
 sky130_fd_sc_hd__mux2_1 _1884_ (.A0(\ram[62][1] ),
    .A1(\ram[63][1] ),
    .S(_0604_),
    .X(_0683_));
 sky130_fd_sc_hd__o221a_1 _1885_ (.A1(_0681_),
    .A2(_0682_),
    .B1(_0683_),
    .B2(_0606_),
    .C1(_0573_),
    .X(_0684_));
 sky130_fd_sc_hd__mux4_1 _1886_ (.A0(\ram[56][1] ),
    .A1(\ram[57][1] ),
    .A2(\ram[58][1] ),
    .A3(\ram[59][1] ),
    .S0(_0608_),
    .S1(_0553_),
    .X(_0685_));
 sky130_fd_sc_hd__and2_1 _1887_ (.A(_0575_),
    .B(_0685_),
    .X(_0686_));
 sky130_fd_sc_hd__o21a_1 _1888_ (.A1(_0684_),
    .A2(_0686_),
    .B1(_0611_),
    .X(_0687_));
 sky130_fd_sc_hd__o31a_1 _1889_ (.A1(_0584_),
    .A2(_0680_),
    .A3(_0687_),
    .B1(_0005_),
    .X(_0688_));
 sky130_fd_sc_hd__mux2_1 _1890_ (.A0(\ram[4][1] ),
    .A1(\ram[5][1] ),
    .S(_0615_),
    .X(_0689_));
 sky130_fd_sc_hd__or2_1 _1891_ (.A(_0614_),
    .B(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__mux2_1 _1892_ (.A0(\ram[6][1] ),
    .A1(\ram[7][1] ),
    .S(_0619_),
    .X(_0691_));
 sky130_fd_sc_hd__o21a_1 _1893_ (.A1(_0618_),
    .A2(_0691_),
    .B1(_0621_),
    .X(_0692_));
 sky130_fd_sc_hd__mux4_1 _1894_ (.A0(\ram[0][1] ),
    .A1(\ram[1][1] ),
    .A2(\ram[2][1] ),
    .A3(\ram[3][1] ),
    .S0(_0623_),
    .S1(_0624_),
    .X(_0693_));
 sky130_fd_sc_hd__a22o_1 _1895_ (.A1(_0690_),
    .A2(_0692_),
    .B1(_0693_),
    .B2(_0626_),
    .X(_0694_));
 sky130_fd_sc_hd__mux2_1 _1896_ (.A0(\ram[20][1] ),
    .A1(\ram[21][1] ),
    .S(_0629_),
    .X(_0695_));
 sky130_fd_sc_hd__or2_1 _1897_ (.A(_0628_),
    .B(_0695_),
    .X(_0696_));
 sky130_fd_sc_hd__mux2_1 _1898_ (.A0(\ram[22][1] ),
    .A1(\ram[23][1] ),
    .S(_0608_),
    .X(_0697_));
 sky130_fd_sc_hd__o21a_1 _1899_ (.A1(_0618_),
    .A2(_0697_),
    .B1(_0544_),
    .X(_0698_));
 sky130_fd_sc_hd__mux4_1 _1900_ (.A0(\ram[16][1] ),
    .A1(\ram[17][1] ),
    .A2(\ram[18][1] ),
    .A3(\ram[19][1] ),
    .S0(_0588_),
    .S1(_0634_),
    .X(_0699_));
 sky130_fd_sc_hd__a22o_1 _1901_ (.A1(_0696_),
    .A2(_0698_),
    .B1(_0699_),
    .B2(_0626_),
    .X(_0700_));
 sky130_fd_sc_hd__mux4_1 _1902_ (.A0(\ram[12][1] ),
    .A1(\ram[13][1] ),
    .A2(\ram[14][1] ),
    .A3(\ram[15][1] ),
    .S0(_0638_),
    .S1(_0624_),
    .X(_0701_));
 sky130_fd_sc_hd__and2b_1 _1903_ (.A_N(_0604_),
    .B(\ram[8][1] ),
    .X(_0702_));
 sky130_fd_sc_hd__a21o_1 _1904_ (.A1(_0641_),
    .A2(\ram[9][1] ),
    .B1(_0550_),
    .X(_0703_));
 sky130_fd_sc_hd__mux2_1 _1905_ (.A0(\ram[10][1] ),
    .A1(\ram[11][1] ),
    .S(_0576_),
    .X(_0704_));
 sky130_fd_sc_hd__o221a_1 _1906_ (.A1(_0702_),
    .A2(_0703_),
    .B1(_0704_),
    .B2(_0644_),
    .C1(_0563_),
    .X(_0705_));
 sky130_fd_sc_hd__a21o_1 _1907_ (.A1(_0637_),
    .A2(_0701_),
    .B1(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__mux4_1 _1908_ (.A0(\ram[28][1] ),
    .A1(\ram[29][1] ),
    .A2(\ram[30][1] ),
    .A3(\ram[31][1] ),
    .S0(_0638_),
    .S1(_0628_),
    .X(_0707_));
 sky130_fd_sc_hd__and2b_1 _1909_ (.A_N(_0649_),
    .B(\ram[24][1] ),
    .X(_0708_));
 sky130_fd_sc_hd__a21o_1 _1910_ (.A1(_0651_),
    .A2(\ram[25][1] ),
    .B1(_0652_),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_1 _1911_ (.A0(\ram[26][1] ),
    .A1(\ram[27][1] ),
    .S(_0619_),
    .X(_0710_));
 sky130_fd_sc_hd__o221a_1 _1912_ (.A1(_0708_),
    .A2(_0709_),
    .B1(_0710_),
    .B2(_0644_),
    .C1(_0645_),
    .X(_0711_));
 sky130_fd_sc_hd__a21o_1 _1913_ (.A1(_0637_),
    .A2(_0707_),
    .B1(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__mux4_2 _1914_ (.A0(_0694_),
    .A1(_0700_),
    .A2(_0706_),
    .A3(_0712_),
    .S0(_0004_),
    .S1(_0543_),
    .X(_0713_));
 sky130_fd_sc_hd__a22o_1 _1915_ (.A1(_0673_),
    .A2(_0688_),
    .B1(_0713_),
    .B2(_0659_),
    .X(net17));
 sky130_fd_sc_hd__mux4_1 _1916_ (.A0(\ram[44][2] ),
    .A1(\ram[45][2] ),
    .A2(\ram[46][2] ),
    .A3(\ram[47][2] ),
    .S0(_0548_),
    .S1(_0551_),
    .X(_0714_));
 sky130_fd_sc_hd__mux2_1 _1917_ (.A0(\ram[40][2] ),
    .A1(\ram[41][2] ),
    .S(_0556_),
    .X(_0715_));
 sky130_fd_sc_hd__or2_1 _1918_ (.A(_0554_),
    .B(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__mux2_1 _1919_ (.A0(\ram[42][2] ),
    .A1(\ram[43][2] ),
    .S(_0561_),
    .X(_0717_));
 sky130_fd_sc_hd__o21a_1 _1920_ (.A1(_0560_),
    .A2(_0717_),
    .B1(_0564_),
    .X(_0718_));
 sky130_fd_sc_hd__a22o_1 _1921_ (.A1(_0546_),
    .A2(_0714_),
    .B1(_0716_),
    .B2(_0718_),
    .X(_0719_));
 sky130_fd_sc_hd__and2b_1 _1922_ (.A_N(_0568_),
    .B(\ram[36][2] ),
    .X(_0720_));
 sky130_fd_sc_hd__a21o_1 _1923_ (.A1(_0602_),
    .A2(\ram[37][2] ),
    .B1(_0570_),
    .X(_0721_));
 sky130_fd_sc_hd__mux2_1 _1924_ (.A0(\ram[38][2] ),
    .A1(\ram[39][2] ),
    .S(_0649_),
    .X(_0722_));
 sky130_fd_sc_hd__o221a_1 _1925_ (.A1(_0720_),
    .A2(_0721_),
    .B1(_0722_),
    .B2(_0606_),
    .C1(_0573_),
    .X(_0723_));
 sky130_fd_sc_hd__mux4_1 _1926_ (.A0(\ram[32][2] ),
    .A1(\ram[33][2] ),
    .A2(\ram[34][2] ),
    .A3(\ram[35][2] ),
    .S0(_0576_),
    .S1(_0577_),
    .X(_0724_));
 sky130_fd_sc_hd__and2_1 _1927_ (.A(_0575_),
    .B(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__o21ba_1 _1928_ (.A1(_0723_),
    .A2(_0725_),
    .B1_N(_0542_),
    .X(_0726_));
 sky130_fd_sc_hd__a211o_1 _1929_ (.A1(_0543_),
    .A2(_0719_),
    .B1(_0726_),
    .C1(_0581_),
    .X(_0727_));
 sky130_fd_sc_hd__buf_4 _1930_ (.A(_0001_),
    .X(_0728_));
 sky130_fd_sc_hd__mux4_1 _1931_ (.A0(\ram[52][2] ),
    .A1(\ram[53][2] ),
    .A2(\ram[54][2] ),
    .A3(\ram[55][2] ),
    .S0(_0547_),
    .S1(_0728_),
    .X(_0729_));
 sky130_fd_sc_hd__and2_1 _1932_ (.A(_0545_),
    .B(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__and2b_1 _1933_ (.A_N(_0588_),
    .B(\ram[48][2] ),
    .X(_0731_));
 sky130_fd_sc_hd__a21o_1 _1934_ (.A1(_0590_),
    .A2(\ram[49][2] ),
    .B1(_0591_),
    .X(_0732_));
 sky130_fd_sc_hd__buf_4 _1935_ (.A(_0555_),
    .X(_0733_));
 sky130_fd_sc_hd__mux2_1 _1936_ (.A0(\ram[50][2] ),
    .A1(\ram[51][2] ),
    .S(_0733_),
    .X(_0734_));
 sky130_fd_sc_hd__o221a_1 _1937_ (.A1(_0731_),
    .A2(_0732_),
    .B1(_0734_),
    .B2(_0595_),
    .C1(_0596_),
    .X(_0735_));
 sky130_fd_sc_hd__o21ba_1 _1938_ (.A1(_0730_),
    .A2(_0735_),
    .B1_N(_0598_),
    .X(_0736_));
 sky130_fd_sc_hd__and2b_1 _1939_ (.A_N(_0600_),
    .B(\ram[60][2] ),
    .X(_0737_));
 sky130_fd_sc_hd__a21o_1 _1940_ (.A1(_0602_),
    .A2(\ram[61][2] ),
    .B1(_0570_),
    .X(_0738_));
 sky130_fd_sc_hd__mux2_1 _1941_ (.A0(\ram[62][2] ),
    .A1(\ram[63][2] ),
    .S(_0604_),
    .X(_0739_));
 sky130_fd_sc_hd__o221a_1 _1942_ (.A1(_0737_),
    .A2(_0738_),
    .B1(_0739_),
    .B2(_0606_),
    .C1(_0585_),
    .X(_0740_));
 sky130_fd_sc_hd__mux4_1 _1943_ (.A0(\ram[56][2] ),
    .A1(\ram[57][2] ),
    .A2(\ram[58][2] ),
    .A3(\ram[59][2] ),
    .S0(_0615_),
    .S1(_0553_),
    .X(_0741_));
 sky130_fd_sc_hd__and2_1 _1944_ (.A(_0596_),
    .B(_0741_),
    .X(_0742_));
 sky130_fd_sc_hd__o21a_1 _1945_ (.A1(_0740_),
    .A2(_0742_),
    .B1(_0542_),
    .X(_0743_));
 sky130_fd_sc_hd__o31a_1 _1946_ (.A1(_0584_),
    .A2(_0736_),
    .A3(_0743_),
    .B1(_0005_),
    .X(_0744_));
 sky130_fd_sc_hd__mux2_1 _1947_ (.A0(\ram[4][2] ),
    .A1(\ram[5][2] ),
    .S(_0615_),
    .X(_0745_));
 sky130_fd_sc_hd__or2_1 _1948_ (.A(_0614_),
    .B(_0745_),
    .X(_0746_));
 sky130_fd_sc_hd__mux2_1 _1949_ (.A0(\ram[6][2] ),
    .A1(\ram[7][2] ),
    .S(_0619_),
    .X(_0747_));
 sky130_fd_sc_hd__o21a_1 _1950_ (.A1(_0618_),
    .A2(_0747_),
    .B1(_0621_),
    .X(_0748_));
 sky130_fd_sc_hd__mux4_1 _1951_ (.A0(\ram[0][2] ),
    .A1(\ram[1][2] ),
    .A2(\ram[2][2] ),
    .A3(\ram[3][2] ),
    .S0(_0623_),
    .S1(_0634_),
    .X(_0749_));
 sky130_fd_sc_hd__a22o_1 _1952_ (.A1(_0746_),
    .A2(_0748_),
    .B1(_0749_),
    .B2(_0626_),
    .X(_0750_));
 sky130_fd_sc_hd__mux2_1 _1953_ (.A0(\ram[20][2] ),
    .A1(\ram[21][2] ),
    .S(_0629_),
    .X(_0751_));
 sky130_fd_sc_hd__or2_1 _1954_ (.A(_0628_),
    .B(_0751_),
    .X(_0752_));
 sky130_fd_sc_hd__mux2_1 _1955_ (.A0(\ram[22][2] ),
    .A1(\ram[23][2] ),
    .S(_0608_),
    .X(_0753_));
 sky130_fd_sc_hd__o21a_1 _1956_ (.A1(_0559_),
    .A2(_0753_),
    .B1(_0544_),
    .X(_0754_));
 sky130_fd_sc_hd__mux4_2 _1957_ (.A0(\ram[16][2] ),
    .A1(\ram[17][2] ),
    .A2(\ram[18][2] ),
    .A3(\ram[19][2] ),
    .S0(_0561_),
    .S1(_0634_),
    .X(_0755_));
 sky130_fd_sc_hd__a22o_1 _1958_ (.A1(_0752_),
    .A2(_0754_),
    .B1(_0755_),
    .B2(_0564_),
    .X(_0756_));
 sky130_fd_sc_hd__mux4_1 _1959_ (.A0(\ram[12][2] ),
    .A1(\ram[13][2] ),
    .A2(\ram[14][2] ),
    .A3(\ram[15][2] ),
    .S0(_0638_),
    .S1(_0624_),
    .X(_0757_));
 sky130_fd_sc_hd__and2b_1 _1960_ (.A_N(_0604_),
    .B(\ram[8][2] ),
    .X(_0758_));
 sky130_fd_sc_hd__a21o_1 _1961_ (.A1(_0641_),
    .A2(\ram[9][2] ),
    .B1(_0550_),
    .X(_0759_));
 sky130_fd_sc_hd__mux2_1 _1962_ (.A0(\ram[10][2] ),
    .A1(\ram[11][2] ),
    .S(_0576_),
    .X(_0760_));
 sky130_fd_sc_hd__o221a_1 _1963_ (.A1(_0758_),
    .A2(_0759_),
    .B1(_0760_),
    .B2(_0644_),
    .C1(_0563_),
    .X(_0761_));
 sky130_fd_sc_hd__a21o_1 _1964_ (.A1(_0637_),
    .A2(_0757_),
    .B1(_0761_),
    .X(_0762_));
 sky130_fd_sc_hd__mux4_1 _1965_ (.A0(\ram[28][2] ),
    .A1(\ram[29][2] ),
    .A2(\ram[30][2] ),
    .A3(\ram[31][2] ),
    .S0(_0638_),
    .S1(_0628_),
    .X(_0763_));
 sky130_fd_sc_hd__and2b_1 _1966_ (.A_N(_0649_),
    .B(\ram[24][2] ),
    .X(_0764_));
 sky130_fd_sc_hd__a21o_1 _1967_ (.A1(_0651_),
    .A2(\ram[25][2] ),
    .B1(_0652_),
    .X(_0765_));
 sky130_fd_sc_hd__mux2_1 _1968_ (.A0(\ram[26][2] ),
    .A1(\ram[27][2] ),
    .S(_0619_),
    .X(_0766_));
 sky130_fd_sc_hd__o221a_1 _1969_ (.A1(_0764_),
    .A2(_0765_),
    .B1(_0766_),
    .B2(_0644_),
    .C1(_0645_),
    .X(_0767_));
 sky130_fd_sc_hd__a21o_1 _1970_ (.A1(_0637_),
    .A2(_0763_),
    .B1(_0767_),
    .X(_0768_));
 sky130_fd_sc_hd__mux4_1 _1971_ (.A0(_0750_),
    .A1(_0756_),
    .A2(_0762_),
    .A3(_0768_),
    .S0(_0004_),
    .S1(_0611_),
    .X(_0769_));
 sky130_fd_sc_hd__a22o_1 _1972_ (.A1(_0727_),
    .A2(_0744_),
    .B1(_0769_),
    .B2(_0659_),
    .X(net18));
 sky130_fd_sc_hd__mux4_1 _1973_ (.A0(\ram[44][3] ),
    .A1(\ram[45][3] ),
    .A2(\ram[46][3] ),
    .A3(\ram[47][3] ),
    .S0(_0548_),
    .S1(_0551_),
    .X(_0770_));
 sky130_fd_sc_hd__mux2_1 _1974_ (.A0(\ram[40][3] ),
    .A1(\ram[41][3] ),
    .S(_0556_),
    .X(_0771_));
 sky130_fd_sc_hd__or2_1 _1975_ (.A(_0554_),
    .B(_0771_),
    .X(_0772_));
 sky130_fd_sc_hd__mux2_1 _1976_ (.A0(\ram[42][3] ),
    .A1(\ram[43][3] ),
    .S(_0561_),
    .X(_0773_));
 sky130_fd_sc_hd__o21a_1 _1977_ (.A1(_0560_),
    .A2(_0773_),
    .B1(_0564_),
    .X(_0774_));
 sky130_fd_sc_hd__a22o_1 _1978_ (.A1(_0546_),
    .A2(_0770_),
    .B1(_0772_),
    .B2(_0774_),
    .X(_0775_));
 sky130_fd_sc_hd__and2b_1 _1979_ (.A_N(_0568_),
    .B(\ram[36][3] ),
    .X(_0776_));
 sky130_fd_sc_hd__a21o_1 _1980_ (.A1(_0602_),
    .A2(\ram[37][3] ),
    .B1(_0570_),
    .X(_0777_));
 sky130_fd_sc_hd__mux2_1 _1981_ (.A0(\ram[38][3] ),
    .A1(\ram[39][3] ),
    .S(_0649_),
    .X(_0778_));
 sky130_fd_sc_hd__o221a_1 _1982_ (.A1(_0776_),
    .A2(_0777_),
    .B1(_0778_),
    .B2(_0606_),
    .C1(_0573_),
    .X(_0779_));
 sky130_fd_sc_hd__mux4_1 _1983_ (.A0(\ram[32][3] ),
    .A1(\ram[33][3] ),
    .A2(\ram[34][3] ),
    .A3(\ram[35][3] ),
    .S0(_0576_),
    .S1(_0577_),
    .X(_0780_));
 sky130_fd_sc_hd__and2_1 _1984_ (.A(_0575_),
    .B(_0780_),
    .X(_0781_));
 sky130_fd_sc_hd__o21ba_1 _1985_ (.A1(_0779_),
    .A2(_0781_),
    .B1_N(_0598_),
    .X(_0782_));
 sky130_fd_sc_hd__a211o_1 _1986_ (.A1(_0543_),
    .A2(_0775_),
    .B1(_0782_),
    .C1(_0581_),
    .X(_0783_));
 sky130_fd_sc_hd__mux4_1 _1987_ (.A0(\ram[52][3] ),
    .A1(\ram[53][3] ),
    .A2(\ram[54][3] ),
    .A3(\ram[55][3] ),
    .S0(_0547_),
    .S1(_0728_),
    .X(_0784_));
 sky130_fd_sc_hd__and2_1 _1988_ (.A(_0545_),
    .B(_0784_),
    .X(_0785_));
 sky130_fd_sc_hd__and2b_1 _1989_ (.A_N(_0588_),
    .B(\ram[48][3] ),
    .X(_0786_));
 sky130_fd_sc_hd__a21o_1 _1990_ (.A1(_0590_),
    .A2(\ram[49][3] ),
    .B1(_0591_),
    .X(_0787_));
 sky130_fd_sc_hd__mux2_1 _1991_ (.A0(\ram[50][3] ),
    .A1(\ram[51][3] ),
    .S(_0733_),
    .X(_0788_));
 sky130_fd_sc_hd__o221a_1 _1992_ (.A1(_0786_),
    .A2(_0787_),
    .B1(_0788_),
    .B2(_0595_),
    .C1(_0596_),
    .X(_0789_));
 sky130_fd_sc_hd__o21ba_1 _1993_ (.A1(_0785_),
    .A2(_0789_),
    .B1_N(_0598_),
    .X(_0790_));
 sky130_fd_sc_hd__and2b_1 _1994_ (.A_N(_0600_),
    .B(\ram[60][3] ),
    .X(_0791_));
 sky130_fd_sc_hd__a21o_1 _1995_ (.A1(_0602_),
    .A2(\ram[61][3] ),
    .B1(_0570_),
    .X(_0792_));
 sky130_fd_sc_hd__mux2_1 _1996_ (.A0(\ram[62][3] ),
    .A1(\ram[63][3] ),
    .S(_0604_),
    .X(_0793_));
 sky130_fd_sc_hd__o221a_1 _1997_ (.A1(_0791_),
    .A2(_0792_),
    .B1(_0793_),
    .B2(_0606_),
    .C1(_0585_),
    .X(_0794_));
 sky130_fd_sc_hd__mux4_1 _1998_ (.A0(\ram[56][3] ),
    .A1(\ram[57][3] ),
    .A2(\ram[58][3] ),
    .A3(\ram[59][3] ),
    .S0(_0615_),
    .S1(_0553_),
    .X(_0795_));
 sky130_fd_sc_hd__and2_1 _1999_ (.A(_0596_),
    .B(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__o21a_1 _2000_ (.A1(_0794_),
    .A2(_0796_),
    .B1(_0542_),
    .X(_0797_));
 sky130_fd_sc_hd__o31a_1 _2001_ (.A1(_0584_),
    .A2(_0790_),
    .A3(_0797_),
    .B1(_0005_),
    .X(_0798_));
 sky130_fd_sc_hd__mux2_1 _2002_ (.A0(\ram[4][3] ),
    .A1(\ram[5][3] ),
    .S(_0615_),
    .X(_0799_));
 sky130_fd_sc_hd__or2_1 _2003_ (.A(_0614_),
    .B(_0799_),
    .X(_0800_));
 sky130_fd_sc_hd__mux2_1 _2004_ (.A0(\ram[6][3] ),
    .A1(\ram[7][3] ),
    .S(_0619_),
    .X(_0801_));
 sky130_fd_sc_hd__o21a_1 _2005_ (.A1(_0618_),
    .A2(_0801_),
    .B1(_0621_),
    .X(_0802_));
 sky130_fd_sc_hd__mux4_1 _2006_ (.A0(\ram[0][3] ),
    .A1(\ram[1][3] ),
    .A2(\ram[2][3] ),
    .A3(\ram[3][3] ),
    .S0(_0623_),
    .S1(_0634_),
    .X(_0803_));
 sky130_fd_sc_hd__a22o_1 _2007_ (.A1(_0800_),
    .A2(_0802_),
    .B1(_0803_),
    .B2(_0626_),
    .X(_0804_));
 sky130_fd_sc_hd__mux2_1 _2008_ (.A0(\ram[20][3] ),
    .A1(\ram[21][3] ),
    .S(_0629_),
    .X(_0805_));
 sky130_fd_sc_hd__or2_1 _2009_ (.A(_0628_),
    .B(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__mux2_1 _2010_ (.A0(\ram[22][3] ),
    .A1(\ram[23][3] ),
    .S(_0608_),
    .X(_0807_));
 sky130_fd_sc_hd__o21a_1 _2011_ (.A1(_0559_),
    .A2(_0807_),
    .B1(_0544_),
    .X(_0808_));
 sky130_fd_sc_hd__mux4_2 _2012_ (.A0(\ram[16][3] ),
    .A1(\ram[17][3] ),
    .A2(\ram[18][3] ),
    .A3(\ram[19][3] ),
    .S0(_0561_),
    .S1(_0634_),
    .X(_0809_));
 sky130_fd_sc_hd__a22o_1 _2013_ (.A1(_0806_),
    .A2(_0808_),
    .B1(_0809_),
    .B2(_0564_),
    .X(_0810_));
 sky130_fd_sc_hd__mux4_1 _2014_ (.A0(\ram[12][3] ),
    .A1(\ram[13][3] ),
    .A2(\ram[14][3] ),
    .A3(\ram[15][3] ),
    .S0(_0600_),
    .S1(_0624_),
    .X(_0811_));
 sky130_fd_sc_hd__and2b_1 _2015_ (.A_N(_0593_),
    .B(\ram[8][3] ),
    .X(_0812_));
 sky130_fd_sc_hd__a21o_1 _2016_ (.A1(_0641_),
    .A2(\ram[9][3] ),
    .B1(_0550_),
    .X(_0813_));
 sky130_fd_sc_hd__mux2_1 _2017_ (.A0(\ram[10][3] ),
    .A1(\ram[11][3] ),
    .S(_0576_),
    .X(_0814_));
 sky130_fd_sc_hd__o221a_1 _2018_ (.A1(_0812_),
    .A2(_0813_),
    .B1(_0814_),
    .B2(_0618_),
    .C1(_0563_),
    .X(_0815_));
 sky130_fd_sc_hd__a21o_1 _2019_ (.A1(_0573_),
    .A2(_0811_),
    .B1(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__mux4_1 _2020_ (.A0(\ram[28][3] ),
    .A1(\ram[29][3] ),
    .A2(\ram[30][3] ),
    .A3(\ram[31][3] ),
    .S0(_0638_),
    .S1(_0624_),
    .X(_0817_));
 sky130_fd_sc_hd__and2b_1 _2021_ (.A_N(_0649_),
    .B(\ram[24][3] ),
    .X(_0818_));
 sky130_fd_sc_hd__a21o_1 _2022_ (.A1(_0651_),
    .A2(\ram[25][3] ),
    .B1(_0652_),
    .X(_0819_));
 sky130_fd_sc_hd__mux2_1 _2023_ (.A0(\ram[26][3] ),
    .A1(\ram[27][3] ),
    .S(_0619_),
    .X(_0820_));
 sky130_fd_sc_hd__o221a_1 _2024_ (.A1(_0818_),
    .A2(_0819_),
    .B1(_0820_),
    .B2(_0644_),
    .C1(_0645_),
    .X(_0821_));
 sky130_fd_sc_hd__a21o_1 _2025_ (.A1(_0637_),
    .A2(_0817_),
    .B1(_0821_),
    .X(_0822_));
 sky130_fd_sc_hd__mux4_2 _2026_ (.A0(_0804_),
    .A1(_0810_),
    .A2(_0816_),
    .A3(_0822_),
    .S0(_0004_),
    .S1(_0611_),
    .X(_0823_));
 sky130_fd_sc_hd__a22o_1 _2027_ (.A1(_0783_),
    .A2(_0798_),
    .B1(_0823_),
    .B2(_0659_),
    .X(net19));
 sky130_fd_sc_hd__mux4_1 _2028_ (.A0(\ram[44][4] ),
    .A1(\ram[45][4] ),
    .A2(\ram[46][4] ),
    .A3(\ram[47][4] ),
    .S0(_0548_),
    .S1(_0551_),
    .X(_0824_));
 sky130_fd_sc_hd__mux2_1 _2029_ (.A0(\ram[40][4] ),
    .A1(\ram[41][4] ),
    .S(_0556_),
    .X(_0825_));
 sky130_fd_sc_hd__or2_1 _2030_ (.A(_0554_),
    .B(_0825_),
    .X(_0826_));
 sky130_fd_sc_hd__mux2_1 _2031_ (.A0(\ram[42][4] ),
    .A1(\ram[43][4] ),
    .S(_0651_),
    .X(_0827_));
 sky130_fd_sc_hd__o21a_1 _2032_ (.A1(_0560_),
    .A2(_0827_),
    .B1(_0564_),
    .X(_0828_));
 sky130_fd_sc_hd__a22o_1 _2033_ (.A1(_0546_),
    .A2(_0824_),
    .B1(_0826_),
    .B2(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__and2b_1 _2034_ (.A_N(_0568_),
    .B(\ram[36][4] ),
    .X(_0830_));
 sky130_fd_sc_hd__a21o_1 _2035_ (.A1(_0602_),
    .A2(\ram[37][4] ),
    .B1(_0570_),
    .X(_0831_));
 sky130_fd_sc_hd__mux2_1 _2036_ (.A0(\ram[38][4] ),
    .A1(\ram[39][4] ),
    .S(_0649_),
    .X(_0832_));
 sky130_fd_sc_hd__o221a_1 _2037_ (.A1(_0830_),
    .A2(_0831_),
    .B1(_0832_),
    .B2(_0606_),
    .C1(_0573_),
    .X(_0833_));
 sky130_fd_sc_hd__mux4_1 _2038_ (.A0(\ram[32][4] ),
    .A1(\ram[33][4] ),
    .A2(\ram[34][4] ),
    .A3(\ram[35][4] ),
    .S0(_0576_),
    .S1(_0553_),
    .X(_0834_));
 sky130_fd_sc_hd__and2_1 _2039_ (.A(_0575_),
    .B(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__o21ba_1 _2040_ (.A1(_0833_),
    .A2(_0835_),
    .B1_N(_0598_),
    .X(_0836_));
 sky130_fd_sc_hd__a211o_1 _2041_ (.A1(_0543_),
    .A2(_0829_),
    .B1(_0836_),
    .C1(_0581_),
    .X(_0837_));
 sky130_fd_sc_hd__mux4_1 _2042_ (.A0(\ram[52][4] ),
    .A1(\ram[53][4] ),
    .A2(\ram[54][4] ),
    .A3(\ram[55][4] ),
    .S0(_0547_),
    .S1(_0728_),
    .X(_0838_));
 sky130_fd_sc_hd__and2_1 _2043_ (.A(_0545_),
    .B(_0838_),
    .X(_0839_));
 sky130_fd_sc_hd__and2b_1 _2044_ (.A_N(_0588_),
    .B(\ram[48][4] ),
    .X(_0840_));
 sky130_fd_sc_hd__a21o_1 _2045_ (.A1(_0568_),
    .A2(\ram[49][4] ),
    .B1(_0591_),
    .X(_0841_));
 sky130_fd_sc_hd__mux2_1 _2046_ (.A0(\ram[50][4] ),
    .A1(\ram[51][4] ),
    .S(_0733_),
    .X(_0842_));
 sky130_fd_sc_hd__o221a_1 _2047_ (.A1(_0840_),
    .A2(_0841_),
    .B1(_0842_),
    .B2(_0595_),
    .C1(_0596_),
    .X(_0843_));
 sky130_fd_sc_hd__o21ba_1 _2048_ (.A1(_0839_),
    .A2(_0843_),
    .B1_N(_0598_),
    .X(_0844_));
 sky130_fd_sc_hd__and2b_1 _2049_ (.A_N(_0600_),
    .B(\ram[60][4] ),
    .X(_0845_));
 sky130_fd_sc_hd__a21o_1 _2050_ (.A1(_0590_),
    .A2(\ram[61][4] ),
    .B1(_0591_),
    .X(_0846_));
 sky130_fd_sc_hd__mux2_1 _2051_ (.A0(\ram[62][4] ),
    .A1(\ram[63][4] ),
    .S(_0604_),
    .X(_0847_));
 sky130_fd_sc_hd__o221a_1 _2052_ (.A1(_0845_),
    .A2(_0846_),
    .B1(_0847_),
    .B2(_0606_),
    .C1(_0585_),
    .X(_0848_));
 sky130_fd_sc_hd__mux4_1 _2053_ (.A0(\ram[56][4] ),
    .A1(\ram[57][4] ),
    .A2(\ram[58][4] ),
    .A3(\ram[59][4] ),
    .S0(_0615_),
    .S1(_0553_),
    .X(_0849_));
 sky130_fd_sc_hd__and2_1 _2054_ (.A(_0596_),
    .B(_0849_),
    .X(_0850_));
 sky130_fd_sc_hd__o21a_1 _2055_ (.A1(_0848_),
    .A2(_0850_),
    .B1(_0542_),
    .X(_0851_));
 sky130_fd_sc_hd__o31a_1 _2056_ (.A1(_0584_),
    .A2(_0844_),
    .A3(_0851_),
    .B1(_0005_),
    .X(_0852_));
 sky130_fd_sc_hd__mux2_1 _2057_ (.A0(\ram[4][4] ),
    .A1(\ram[5][4] ),
    .S(_0615_),
    .X(_0853_));
 sky130_fd_sc_hd__or2_1 _2058_ (.A(_0614_),
    .B(_0853_),
    .X(_0854_));
 sky130_fd_sc_hd__mux2_1 _2059_ (.A0(\ram[6][4] ),
    .A1(\ram[7][4] ),
    .S(_0619_),
    .X(_0855_));
 sky130_fd_sc_hd__o21a_1 _2060_ (.A1(_0618_),
    .A2(_0855_),
    .B1(_0621_),
    .X(_0856_));
 sky130_fd_sc_hd__mux4_1 _2061_ (.A0(\ram[0][4] ),
    .A1(\ram[1][4] ),
    .A2(\ram[2][4] ),
    .A3(\ram[3][4] ),
    .S0(_0623_),
    .S1(_0634_),
    .X(_0857_));
 sky130_fd_sc_hd__a22o_1 _2062_ (.A1(_0854_),
    .A2(_0856_),
    .B1(_0857_),
    .B2(_0626_),
    .X(_0858_));
 sky130_fd_sc_hd__mux2_1 _2063_ (.A0(\ram[20][4] ),
    .A1(\ram[21][4] ),
    .S(_0629_),
    .X(_0859_));
 sky130_fd_sc_hd__or2_1 _2064_ (.A(_0628_),
    .B(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__mux2_1 _2065_ (.A0(\ram[22][4] ),
    .A1(\ram[23][4] ),
    .S(_0608_),
    .X(_0861_));
 sky130_fd_sc_hd__o21a_1 _2066_ (.A1(_0559_),
    .A2(_0861_),
    .B1(_0544_),
    .X(_0862_));
 sky130_fd_sc_hd__mux4_2 _2067_ (.A0(\ram[16][4] ),
    .A1(\ram[17][4] ),
    .A2(\ram[18][4] ),
    .A3(\ram[19][4] ),
    .S0(_0561_),
    .S1(_0634_),
    .X(_0863_));
 sky130_fd_sc_hd__a22o_1 _2068_ (.A1(_0860_),
    .A2(_0862_),
    .B1(_0863_),
    .B2(_0564_),
    .X(_0864_));
 sky130_fd_sc_hd__mux4_1 _2069_ (.A0(\ram[12][4] ),
    .A1(\ram[13][4] ),
    .A2(\ram[14][4] ),
    .A3(\ram[15][4] ),
    .S0(_0600_),
    .S1(_0624_),
    .X(_0865_));
 sky130_fd_sc_hd__and2b_1 _2070_ (.A_N(_0593_),
    .B(\ram[8][4] ),
    .X(_0866_));
 sky130_fd_sc_hd__a21o_1 _2071_ (.A1(_0641_),
    .A2(\ram[9][4] ),
    .B1(_0550_),
    .X(_0867_));
 sky130_fd_sc_hd__mux2_1 _2072_ (.A0(\ram[10][4] ),
    .A1(\ram[11][4] ),
    .S(_0576_),
    .X(_0868_));
 sky130_fd_sc_hd__o221a_1 _2073_ (.A1(_0866_),
    .A2(_0867_),
    .B1(_0868_),
    .B2(_0618_),
    .C1(_0563_),
    .X(_0869_));
 sky130_fd_sc_hd__a21o_1 _2074_ (.A1(_0573_),
    .A2(_0865_),
    .B1(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__mux4_1 _2075_ (.A0(\ram[28][4] ),
    .A1(\ram[29][4] ),
    .A2(\ram[30][4] ),
    .A3(\ram[31][4] ),
    .S0(_0638_),
    .S1(_0624_),
    .X(_0871_));
 sky130_fd_sc_hd__and2b_1 _2076_ (.A_N(_0649_),
    .B(\ram[24][4] ),
    .X(_0872_));
 sky130_fd_sc_hd__a21o_1 _2077_ (.A1(_0651_),
    .A2(\ram[25][4] ),
    .B1(_0652_),
    .X(_0873_));
 sky130_fd_sc_hd__mux2_1 _2078_ (.A0(\ram[26][4] ),
    .A1(\ram[27][4] ),
    .S(_0619_),
    .X(_0874_));
 sky130_fd_sc_hd__o221a_1 _2079_ (.A1(_0872_),
    .A2(_0873_),
    .B1(_0874_),
    .B2(_0644_),
    .C1(_0645_),
    .X(_0875_));
 sky130_fd_sc_hd__a21o_1 _2080_ (.A1(_0637_),
    .A2(_0871_),
    .B1(_0875_),
    .X(_0876_));
 sky130_fd_sc_hd__mux4_1 _2081_ (.A0(_0858_),
    .A1(_0864_),
    .A2(_0870_),
    .A3(_0876_),
    .S0(_0004_),
    .S1(_0611_),
    .X(_0877_));
 sky130_fd_sc_hd__a22o_1 _2082_ (.A1(_0837_),
    .A2(_0852_),
    .B1(_0877_),
    .B2(_0659_),
    .X(net20));
 sky130_fd_sc_hd__mux4_1 _2083_ (.A0(\ram[44][5] ),
    .A1(\ram[45][5] ),
    .A2(\ram[46][5] ),
    .A3(\ram[47][5] ),
    .S0(_0548_),
    .S1(_0551_),
    .X(_0878_));
 sky130_fd_sc_hd__mux2_1 _2084_ (.A0(\ram[40][5] ),
    .A1(\ram[41][5] ),
    .S(_0556_),
    .X(_0879_));
 sky130_fd_sc_hd__or2_1 _2085_ (.A(_0554_),
    .B(_0879_),
    .X(_0880_));
 sky130_fd_sc_hd__mux2_1 _2086_ (.A0(\ram[42][5] ),
    .A1(\ram[43][5] ),
    .S(_0651_),
    .X(_0881_));
 sky130_fd_sc_hd__o21a_1 _2087_ (.A1(_0560_),
    .A2(_0881_),
    .B1(_0564_),
    .X(_0882_));
 sky130_fd_sc_hd__a22o_1 _2088_ (.A1(_0546_),
    .A2(_0878_),
    .B1(_0880_),
    .B2(_0882_),
    .X(_0883_));
 sky130_fd_sc_hd__and2b_1 _2089_ (.A_N(_0568_),
    .B(\ram[36][5] ),
    .X(_0884_));
 sky130_fd_sc_hd__a21o_1 _2090_ (.A1(_0602_),
    .A2(\ram[37][5] ),
    .B1(_0570_),
    .X(_0885_));
 sky130_fd_sc_hd__mux2_1 _2091_ (.A0(\ram[38][5] ),
    .A1(\ram[39][5] ),
    .S(_0649_),
    .X(_0886_));
 sky130_fd_sc_hd__o221a_1 _2092_ (.A1(_0884_),
    .A2(_0885_),
    .B1(_0886_),
    .B2(_0606_),
    .C1(_0573_),
    .X(_0887_));
 sky130_fd_sc_hd__mux4_1 _2093_ (.A0(\ram[32][5] ),
    .A1(\ram[33][5] ),
    .A2(\ram[34][5] ),
    .A3(\ram[35][5] ),
    .S0(_0608_),
    .S1(_0553_),
    .X(_0888_));
 sky130_fd_sc_hd__and2_1 _2094_ (.A(_0575_),
    .B(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__o21ba_1 _2095_ (.A1(_0887_),
    .A2(_0889_),
    .B1_N(_0598_),
    .X(_0890_));
 sky130_fd_sc_hd__a211o_1 _2096_ (.A1(_0543_),
    .A2(_0883_),
    .B1(_0890_),
    .C1(_0581_),
    .X(_0891_));
 sky130_fd_sc_hd__mux4_1 _2097_ (.A0(\ram[52][5] ),
    .A1(\ram[53][5] ),
    .A2(\ram[54][5] ),
    .A3(\ram[55][5] ),
    .S0(_0547_),
    .S1(_0728_),
    .X(_0892_));
 sky130_fd_sc_hd__and2_1 _2098_ (.A(_0545_),
    .B(_0892_),
    .X(_0893_));
 sky130_fd_sc_hd__and2b_1 _2099_ (.A_N(_0588_),
    .B(\ram[48][5] ),
    .X(_0894_));
 sky130_fd_sc_hd__a21o_1 _2100_ (.A1(_0568_),
    .A2(\ram[49][5] ),
    .B1(_0591_),
    .X(_0895_));
 sky130_fd_sc_hd__mux2_1 _2101_ (.A0(\ram[50][5] ),
    .A1(\ram[51][5] ),
    .S(_0733_),
    .X(_0896_));
 sky130_fd_sc_hd__o221a_1 _2102_ (.A1(_0894_),
    .A2(_0895_),
    .B1(_0896_),
    .B2(_0595_),
    .C1(_0596_),
    .X(_0897_));
 sky130_fd_sc_hd__o21ba_1 _2103_ (.A1(_0893_),
    .A2(_0897_),
    .B1_N(_0003_),
    .X(_0898_));
 sky130_fd_sc_hd__and2b_1 _2104_ (.A_N(_0600_),
    .B(\ram[60][5] ),
    .X(_0899_));
 sky130_fd_sc_hd__a21o_1 _2105_ (.A1(_0590_),
    .A2(\ram[61][5] ),
    .B1(_0591_),
    .X(_0900_));
 sky130_fd_sc_hd__mux2_1 _2106_ (.A0(\ram[62][5] ),
    .A1(\ram[63][5] ),
    .S(_0604_),
    .X(_0901_));
 sky130_fd_sc_hd__o221a_1 _2107_ (.A1(_0899_),
    .A2(_0900_),
    .B1(_0901_),
    .B2(_0606_),
    .C1(_0585_),
    .X(_0902_));
 sky130_fd_sc_hd__mux4_1 _2108_ (.A0(\ram[56][5] ),
    .A1(\ram[57][5] ),
    .A2(\ram[58][5] ),
    .A3(\ram[59][5] ),
    .S0(_0615_),
    .S1(_0652_),
    .X(_0903_));
 sky130_fd_sc_hd__and2_1 _2109_ (.A(_0596_),
    .B(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__o21a_1 _2110_ (.A1(_0902_),
    .A2(_0904_),
    .B1(_0542_),
    .X(_0905_));
 sky130_fd_sc_hd__o31a_1 _2111_ (.A1(_0584_),
    .A2(_0898_),
    .A3(_0905_),
    .B1(_0005_),
    .X(_0906_));
 sky130_fd_sc_hd__mux4_1 _2112_ (.A0(\ram[20][5] ),
    .A1(\ram[21][5] ),
    .A2(\ram[22][5] ),
    .A3(\ram[23][5] ),
    .S0(_0638_),
    .S1(_0628_),
    .X(_0907_));
 sky130_fd_sc_hd__and2b_1 _2113_ (.A_N(_0649_),
    .B(\ram[16][5] ),
    .X(_0908_));
 sky130_fd_sc_hd__a21o_1 _2114_ (.A1(_0651_),
    .A2(\ram[17][5] ),
    .B1(_0652_),
    .X(_0909_));
 sky130_fd_sc_hd__mux2_1 _2115_ (.A0(\ram[18][5] ),
    .A1(\ram[19][5] ),
    .S(_0654_),
    .X(_0910_));
 sky130_fd_sc_hd__o221a_1 _2116_ (.A1(_0908_),
    .A2(_0909_),
    .B1(_0910_),
    .B2(_0644_),
    .C1(_0645_),
    .X(_0911_));
 sky130_fd_sc_hd__a21o_1 _2117_ (.A1(_0637_),
    .A2(_0907_),
    .B1(_0911_),
    .X(_0912_));
 sky130_fd_sc_hd__mux2_1 _2118_ (.A0(\ram[28][5] ),
    .A1(\ram[29][5] ),
    .S(_0629_),
    .X(_0913_));
 sky130_fd_sc_hd__or2_1 _2119_ (.A(_0628_),
    .B(_0913_),
    .X(_0914_));
 sky130_fd_sc_hd__mux2_1 _2120_ (.A0(\ram[30][5] ),
    .A1(\ram[31][5] ),
    .S(_0608_),
    .X(_0915_));
 sky130_fd_sc_hd__o21a_1 _2121_ (.A1(_0559_),
    .A2(_0915_),
    .B1(_0544_),
    .X(_0916_));
 sky130_fd_sc_hd__mux4_1 _2122_ (.A0(\ram[24][5] ),
    .A1(\ram[25][5] ),
    .A2(\ram[26][5] ),
    .A3(\ram[27][5] ),
    .S0(_0561_),
    .S1(_0634_),
    .X(_0917_));
 sky130_fd_sc_hd__a22o_1 _2123_ (.A1(_0914_),
    .A2(_0916_),
    .B1(_0917_),
    .B2(_0564_),
    .X(_0918_));
 sky130_fd_sc_hd__mux2_1 _2124_ (.A0(\ram[4][5] ),
    .A1(\ram[5][5] ),
    .S(_0615_),
    .X(_0919_));
 sky130_fd_sc_hd__or2_1 _2125_ (.A(_0614_),
    .B(_0919_),
    .X(_0920_));
 sky130_fd_sc_hd__mux2_1 _2126_ (.A0(\ram[6][5] ),
    .A1(\ram[7][5] ),
    .S(_0608_),
    .X(_0921_));
 sky130_fd_sc_hd__o21a_1 _2127_ (.A1(_0618_),
    .A2(_0921_),
    .B1(_0621_),
    .X(_0922_));
 sky130_fd_sc_hd__mux4_1 _2128_ (.A0(\ram[0][5] ),
    .A1(\ram[1][5] ),
    .A2(\ram[2][5] ),
    .A3(\ram[3][5] ),
    .S0(_0623_),
    .S1(_0634_),
    .X(_0923_));
 sky130_fd_sc_hd__a22o_1 _2129_ (.A1(_0920_),
    .A2(_0922_),
    .B1(_0923_),
    .B2(_0626_),
    .X(_0924_));
 sky130_fd_sc_hd__mux4_1 _2130_ (.A0(\ram[12][5] ),
    .A1(\ram[13][5] ),
    .A2(\ram[14][5] ),
    .A3(\ram[15][5] ),
    .S0(_0638_),
    .S1(_0624_),
    .X(_0925_));
 sky130_fd_sc_hd__and2b_1 _2131_ (.A_N(_0604_),
    .B(\ram[8][5] ),
    .X(_0926_));
 sky130_fd_sc_hd__a21o_1 _2132_ (.A1(_0641_),
    .A2(\ram[9][5] ),
    .B1(_0652_),
    .X(_0927_));
 sky130_fd_sc_hd__mux2_1 _2133_ (.A0(\ram[10][5] ),
    .A1(\ram[11][5] ),
    .S(_0619_),
    .X(_0928_));
 sky130_fd_sc_hd__o221a_1 _2134_ (.A1(_0926_),
    .A2(_0927_),
    .B1(_0928_),
    .B2(_0644_),
    .C1(_0645_),
    .X(_0929_));
 sky130_fd_sc_hd__a21o_1 _2135_ (.A1(_0637_),
    .A2(_0925_),
    .B1(_0929_),
    .X(_0930_));
 sky130_fd_sc_hd__mux4_1 _2136_ (.A0(_0912_),
    .A1(_0918_),
    .A2(_0924_),
    .A3(_0930_),
    .S0(_0611_),
    .S1(_0584_),
    .X(_0931_));
 sky130_fd_sc_hd__a22o_1 _2137_ (.A1(_0891_),
    .A2(_0906_),
    .B1(_0931_),
    .B2(_0659_),
    .X(net21));
 sky130_fd_sc_hd__mux2_1 _2138_ (.A0(\ram[28][6] ),
    .A1(\ram[29][6] ),
    .S(_0654_),
    .X(_0932_));
 sky130_fd_sc_hd__or2_1 _2139_ (.A(_0551_),
    .B(_0932_),
    .X(_0933_));
 sky130_fd_sc_hd__clkbuf_4 _2140_ (.A(_0559_),
    .X(_0934_));
 sky130_fd_sc_hd__mux2_1 _2141_ (.A0(\ram[30][6] ),
    .A1(\ram[31][6] ),
    .S(_0654_),
    .X(_0935_));
 sky130_fd_sc_hd__o21a_1 _2142_ (.A1(_0934_),
    .A2(_0935_),
    .B1(_0621_),
    .X(_0936_));
 sky130_fd_sc_hd__mux4_1 _2143_ (.A0(\ram[24][6] ),
    .A1(\ram[25][6] ),
    .A2(\ram[26][6] ),
    .A3(\ram[27][6] ),
    .S0(_0602_),
    .S1(_0614_),
    .X(_0937_));
 sky130_fd_sc_hd__a22o_1 _2144_ (.A1(_0933_),
    .A2(_0936_),
    .B1(_0937_),
    .B2(_0626_),
    .X(_0938_));
 sky130_fd_sc_hd__mux4_1 _2145_ (.A0(\ram[20][6] ),
    .A1(\ram[21][6] ),
    .A2(\ram[22][6] ),
    .A3(\ram[23][6] ),
    .S0(_0567_),
    .S1(_0728_),
    .X(_0939_));
 sky130_fd_sc_hd__and2_1 _2146_ (.A(_0621_),
    .B(_0939_),
    .X(_0940_));
 sky130_fd_sc_hd__and2b_1 _2147_ (.A_N(_0641_),
    .B(\ram[16][6] ),
    .X(_0941_));
 sky130_fd_sc_hd__a21o_1 _2148_ (.A1(_0588_),
    .A2(\ram[17][6] ),
    .B1(_0553_),
    .X(_0942_));
 sky130_fd_sc_hd__mux2_1 _2149_ (.A0(\ram[18][6] ),
    .A1(\ram[19][6] ),
    .S(_0654_),
    .X(_0943_));
 sky130_fd_sc_hd__clkbuf_4 _2150_ (.A(_0563_),
    .X(_0944_));
 sky130_fd_sc_hd__o221a_1 _2151_ (.A1(_0941_),
    .A2(_0942_),
    .B1(_0943_),
    .B2(_0934_),
    .C1(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__o21ba_1 _2152_ (.A1(_0940_),
    .A2(_0945_),
    .B1_N(_0003_),
    .X(_0946_));
 sky130_fd_sc_hd__a211o_1 _2153_ (.A1(_0611_),
    .A2(_0938_),
    .B1(_0946_),
    .C1(_0584_),
    .X(_0947_));
 sky130_fd_sc_hd__mux4_1 _2154_ (.A0(\ram[12][6] ),
    .A1(\ram[13][6] ),
    .A2(\ram[14][6] ),
    .A3(\ram[15][6] ),
    .S0(_0590_),
    .S1(_0614_),
    .X(_0948_));
 sky130_fd_sc_hd__mux2_1 _2155_ (.A0(\ram[8][6] ),
    .A1(\ram[9][6] ),
    .S(_0733_),
    .X(_0949_));
 sky130_fd_sc_hd__or2_1 _2156_ (.A(_0554_),
    .B(_0949_),
    .X(_0950_));
 sky130_fd_sc_hd__mux2_1 _2157_ (.A0(\ram[10][6] ),
    .A1(\ram[11][6] ),
    .S(_0593_),
    .X(_0951_));
 sky130_fd_sc_hd__o21a_1 _2158_ (.A1(_0595_),
    .A2(_0951_),
    .B1(_0944_),
    .X(_0952_));
 sky130_fd_sc_hd__a22o_1 _2159_ (.A1(_0546_),
    .A2(_0948_),
    .B1(_0950_),
    .B2(_0952_),
    .X(_0953_));
 sky130_fd_sc_hd__and2b_1 _2160_ (.A_N(_0641_),
    .B(\ram[4][6] ),
    .X(_0954_));
 sky130_fd_sc_hd__a21o_1 _2161_ (.A1(_0623_),
    .A2(\ram[5][6] ),
    .B1(_0577_),
    .X(_0955_));
 sky130_fd_sc_hd__mux2_1 _2162_ (.A0(\ram[6][6] ),
    .A1(\ram[7][6] ),
    .S(_0654_),
    .X(_0956_));
 sky130_fd_sc_hd__o221a_1 _2163_ (.A1(_0954_),
    .A2(_0955_),
    .B1(_0956_),
    .B2(_0934_),
    .C1(_0545_),
    .X(_0957_));
 sky130_fd_sc_hd__mux4_1 _2164_ (.A0(\ram[0][6] ),
    .A1(\ram[1][6] ),
    .A2(\ram[2][6] ),
    .A3(\ram[3][6] ),
    .S0(_0547_),
    .S1(_0728_),
    .X(_0958_));
 sky130_fd_sc_hd__and2_1 _2165_ (.A(_0645_),
    .B(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__o21ba_1 _2166_ (.A1(_0957_),
    .A2(_0959_),
    .B1_N(_0003_),
    .X(_0960_));
 sky130_fd_sc_hd__a211o_1 _2167_ (.A1(_0611_),
    .A2(_0953_),
    .B1(_0960_),
    .C1(_0581_),
    .X(_0961_));
 sky130_fd_sc_hd__mux4_1 _2168_ (.A0(\ram[60][6] ),
    .A1(\ram[61][6] ),
    .A2(\ram[62][6] ),
    .A3(\ram[63][6] ),
    .S0(_0548_),
    .S1(_0551_),
    .X(_0962_));
 sky130_fd_sc_hd__mux2_1 _2169_ (.A0(\ram[56][6] ),
    .A1(\ram[57][6] ),
    .S(_0593_),
    .X(_0963_));
 sky130_fd_sc_hd__or2_1 _2170_ (.A(_0554_),
    .B(_0963_),
    .X(_0964_));
 sky130_fd_sc_hd__mux2_1 _2171_ (.A0(\ram[58][6] ),
    .A1(\ram[59][6] ),
    .S(_0556_),
    .X(_0965_));
 sky130_fd_sc_hd__o21a_1 _2172_ (.A1(_0560_),
    .A2(_0965_),
    .B1(_0575_),
    .X(_0966_));
 sky130_fd_sc_hd__a22o_1 _2173_ (.A1(_0546_),
    .A2(_0962_),
    .B1(_0964_),
    .B2(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__and2b_1 _2174_ (.A_N(_0623_),
    .B(\ram[52][6] ),
    .X(_0968_));
 sky130_fd_sc_hd__a21o_1 _2175_ (.A1(_0590_),
    .A2(\ram[53][6] ),
    .B1(_0591_),
    .X(_0969_));
 sky130_fd_sc_hd__mux2_1 _2176_ (.A0(\ram[54][6] ),
    .A1(\ram[55][6] ),
    .S(_0593_),
    .X(_0970_));
 sky130_fd_sc_hd__o221a_1 _2177_ (.A1(_0968_),
    .A2(_0969_),
    .B1(_0970_),
    .B2(_0595_),
    .C1(_0585_),
    .X(_0971_));
 sky130_fd_sc_hd__mux4_1 _2178_ (.A0(\ram[48][6] ),
    .A1(\ram[49][6] ),
    .A2(\ram[50][6] ),
    .A3(\ram[51][6] ),
    .S0(_0629_),
    .S1(_0652_),
    .X(_0972_));
 sky130_fd_sc_hd__and2_1 _2179_ (.A(_0944_),
    .B(_0972_),
    .X(_0973_));
 sky130_fd_sc_hd__o21ba_1 _2180_ (.A1(_0971_),
    .A2(_0973_),
    .B1_N(_0598_),
    .X(_0974_));
 sky130_fd_sc_hd__a211o_1 _2181_ (.A1(_0543_),
    .A2(_0967_),
    .B1(_0974_),
    .C1(_0584_),
    .X(_0975_));
 sky130_fd_sc_hd__mux4_1 _2182_ (.A0(\ram[44][6] ),
    .A1(\ram[45][6] ),
    .A2(\ram[46][6] ),
    .A3(\ram[47][6] ),
    .S0(_0567_),
    .S1(_0728_),
    .X(_0976_));
 sky130_fd_sc_hd__and2_1 _2183_ (.A(_0545_),
    .B(_0976_),
    .X(_0977_));
 sky130_fd_sc_hd__and2b_1 _2184_ (.A_N(_0651_),
    .B(\ram[40][6] ),
    .X(_0978_));
 sky130_fd_sc_hd__a21o_1 _2185_ (.A1(_0600_),
    .A2(\ram[41][6] ),
    .B1(_0577_),
    .X(_0979_));
 sky130_fd_sc_hd__mux2_1 _2186_ (.A0(\ram[42][6] ),
    .A1(\ram[43][6] ),
    .S(_0733_),
    .X(_0980_));
 sky130_fd_sc_hd__o221a_1 _2187_ (.A1(_0978_),
    .A2(_0979_),
    .B1(_0980_),
    .B2(_0934_),
    .C1(_0944_),
    .X(_0981_));
 sky130_fd_sc_hd__o21a_1 _2188_ (.A1(_0977_),
    .A2(_0981_),
    .B1(_0542_),
    .X(_0982_));
 sky130_fd_sc_hd__and2b_1 _2189_ (.A_N(_0561_),
    .B(\ram[36][6] ),
    .X(_0983_));
 sky130_fd_sc_hd__a21o_1 _2190_ (.A1(_0568_),
    .A2(\ram[37][6] ),
    .B1(_0577_),
    .X(_0984_));
 sky130_fd_sc_hd__mux2_1 _2191_ (.A0(\ram[38][6] ),
    .A1(\ram[39][6] ),
    .S(_0733_),
    .X(_0985_));
 sky130_fd_sc_hd__o221a_1 _2192_ (.A1(_0983_),
    .A2(_0984_),
    .B1(_0985_),
    .B2(_0934_),
    .C1(_0585_),
    .X(_0986_));
 sky130_fd_sc_hd__mux4_1 _2193_ (.A0(\ram[32][6] ),
    .A1(\ram[33][6] ),
    .A2(\ram[34][6] ),
    .A3(\ram[35][6] ),
    .S0(_0629_),
    .S1(_0550_),
    .X(_0987_));
 sky130_fd_sc_hd__and2_1 _2194_ (.A(_0944_),
    .B(_0987_),
    .X(_0988_));
 sky130_fd_sc_hd__o21ba_1 _2195_ (.A1(_0986_),
    .A2(_0988_),
    .B1_N(_0003_),
    .X(_0989_));
 sky130_fd_sc_hd__o31a_1 _2196_ (.A1(_0581_),
    .A2(_0982_),
    .A3(_0989_),
    .B1(_0005_),
    .X(_0990_));
 sky130_fd_sc_hd__a32o_1 _2197_ (.A1(_0659_),
    .A2(_0947_),
    .A3(_0961_),
    .B1(_0975_),
    .B2(_0990_),
    .X(net22));
 sky130_fd_sc_hd__mux2_1 _2198_ (.A0(\ram[28][7] ),
    .A1(\ram[29][7] ),
    .S(_0654_),
    .X(_0991_));
 sky130_fd_sc_hd__or2_1 _2199_ (.A(_0551_),
    .B(_0991_),
    .X(_0992_));
 sky130_fd_sc_hd__mux2_1 _2200_ (.A0(\ram[30][7] ),
    .A1(\ram[31][7] ),
    .S(_0654_),
    .X(_0993_));
 sky130_fd_sc_hd__o21a_1 _2201_ (.A1(_0934_),
    .A2(_0993_),
    .B1(_0621_),
    .X(_0994_));
 sky130_fd_sc_hd__mux4_1 _2202_ (.A0(\ram[24][7] ),
    .A1(\ram[25][7] ),
    .A2(\ram[26][7] ),
    .A3(\ram[27][7] ),
    .S0(_0602_),
    .S1(_0614_),
    .X(_0995_));
 sky130_fd_sc_hd__a22o_1 _2203_ (.A1(_0992_),
    .A2(_0994_),
    .B1(_0995_),
    .B2(_0626_),
    .X(_0996_));
 sky130_fd_sc_hd__mux4_1 _2204_ (.A0(\ram[20][7] ),
    .A1(\ram[21][7] ),
    .A2(\ram[22][7] ),
    .A3(\ram[23][7] ),
    .S0(_0567_),
    .S1(_0728_),
    .X(_0997_));
 sky130_fd_sc_hd__and2_1 _2205_ (.A(_0621_),
    .B(_0997_),
    .X(_0998_));
 sky130_fd_sc_hd__and2b_1 _2206_ (.A_N(_0641_),
    .B(\ram[16][7] ),
    .X(_0999_));
 sky130_fd_sc_hd__a21o_1 _2207_ (.A1(_0588_),
    .A2(\ram[17][7] ),
    .B1(_0553_),
    .X(_1000_));
 sky130_fd_sc_hd__mux2_1 _2208_ (.A0(\ram[18][7] ),
    .A1(\ram[19][7] ),
    .S(_0654_),
    .X(_1001_));
 sky130_fd_sc_hd__o221a_1 _2209_ (.A1(_0999_),
    .A2(_1000_),
    .B1(_1001_),
    .B2(_0934_),
    .C1(_0944_),
    .X(_1002_));
 sky130_fd_sc_hd__o21ba_1 _2210_ (.A1(_0998_),
    .A2(_1002_),
    .B1_N(_0003_),
    .X(_1003_));
 sky130_fd_sc_hd__a211o_1 _2211_ (.A1(_0611_),
    .A2(_0996_),
    .B1(_1003_),
    .C1(_0583_),
    .X(_1004_));
 sky130_fd_sc_hd__mux4_1 _2212_ (.A0(\ram[12][7] ),
    .A1(\ram[13][7] ),
    .A2(\ram[14][7] ),
    .A3(\ram[15][7] ),
    .S0(_0590_),
    .S1(_0614_),
    .X(_1005_));
 sky130_fd_sc_hd__mux2_1 _2213_ (.A0(\ram[8][7] ),
    .A1(\ram[9][7] ),
    .S(_0733_),
    .X(_1006_));
 sky130_fd_sc_hd__or2_1 _2214_ (.A(_0554_),
    .B(_1006_),
    .X(_1007_));
 sky130_fd_sc_hd__mux2_1 _2215_ (.A0(\ram[10][7] ),
    .A1(\ram[11][7] ),
    .S(_0593_),
    .X(_1008_));
 sky130_fd_sc_hd__o21a_1 _2216_ (.A1(_0595_),
    .A2(_1008_),
    .B1(_0944_),
    .X(_1009_));
 sky130_fd_sc_hd__a22o_1 _2217_ (.A1(_0546_),
    .A2(_1005_),
    .B1(_1007_),
    .B2(_1009_),
    .X(_1010_));
 sky130_fd_sc_hd__and2b_1 _2218_ (.A_N(_0641_),
    .B(\ram[4][7] ),
    .X(_1011_));
 sky130_fd_sc_hd__a21o_1 _2219_ (.A1(_0623_),
    .A2(\ram[5][7] ),
    .B1(_0577_),
    .X(_1012_));
 sky130_fd_sc_hd__mux2_1 _2220_ (.A0(\ram[6][7] ),
    .A1(\ram[7][7] ),
    .S(_0654_),
    .X(_1013_));
 sky130_fd_sc_hd__o221a_1 _2221_ (.A1(_1011_),
    .A2(_1012_),
    .B1(_1013_),
    .B2(_0934_),
    .C1(_0545_),
    .X(_1014_));
 sky130_fd_sc_hd__mux4_1 _2222_ (.A0(\ram[0][7] ),
    .A1(\ram[1][7] ),
    .A2(\ram[2][7] ),
    .A3(\ram[3][7] ),
    .S0(_0547_),
    .S1(_0728_),
    .X(_1015_));
 sky130_fd_sc_hd__and2_1 _2223_ (.A(_0645_),
    .B(_1015_),
    .X(_1016_));
 sky130_fd_sc_hd__o21ba_1 _2224_ (.A1(_1014_),
    .A2(_1016_),
    .B1_N(_0003_),
    .X(_1017_));
 sky130_fd_sc_hd__a211o_1 _2225_ (.A1(_0611_),
    .A2(_1010_),
    .B1(_1017_),
    .C1(_0581_),
    .X(_1018_));
 sky130_fd_sc_hd__mux4_1 _2226_ (.A0(\ram[60][7] ),
    .A1(\ram[61][7] ),
    .A2(\ram[62][7] ),
    .A3(\ram[63][7] ),
    .S0(_0548_),
    .S1(_0551_),
    .X(_1019_));
 sky130_fd_sc_hd__mux2_1 _2227_ (.A0(\ram[56][7] ),
    .A1(\ram[57][7] ),
    .S(_0593_),
    .X(_1020_));
 sky130_fd_sc_hd__or2_1 _2228_ (.A(_0554_),
    .B(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__mux2_1 _2229_ (.A0(\ram[58][7] ),
    .A1(\ram[59][7] ),
    .S(_0556_),
    .X(_1022_));
 sky130_fd_sc_hd__o21a_1 _2230_ (.A1(_0560_),
    .A2(_1022_),
    .B1(_0575_),
    .X(_1023_));
 sky130_fd_sc_hd__a22o_1 _2231_ (.A1(_0546_),
    .A2(_1019_),
    .B1(_1021_),
    .B2(_1023_),
    .X(_1024_));
 sky130_fd_sc_hd__and2b_1 _2232_ (.A_N(_0623_),
    .B(\ram[52][7] ),
    .X(_1025_));
 sky130_fd_sc_hd__a21o_1 _2233_ (.A1(_0590_),
    .A2(\ram[53][7] ),
    .B1(_0591_),
    .X(_1026_));
 sky130_fd_sc_hd__mux2_1 _2234_ (.A0(\ram[54][7] ),
    .A1(\ram[55][7] ),
    .S(_0593_),
    .X(_1027_));
 sky130_fd_sc_hd__o221a_1 _2235_ (.A1(_1025_),
    .A2(_1026_),
    .B1(_1027_),
    .B2(_0595_),
    .C1(_0585_),
    .X(_1028_));
 sky130_fd_sc_hd__mux4_1 _2236_ (.A0(\ram[48][7] ),
    .A1(\ram[49][7] ),
    .A2(\ram[50][7] ),
    .A3(\ram[51][7] ),
    .S0(_0629_),
    .S1(_0652_),
    .X(_1029_));
 sky130_fd_sc_hd__and2_1 _2237_ (.A(_0944_),
    .B(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__o21ba_1 _2238_ (.A1(_1028_),
    .A2(_1030_),
    .B1_N(_0598_),
    .X(_1031_));
 sky130_fd_sc_hd__a211o_1 _2239_ (.A1(_0543_),
    .A2(_1024_),
    .B1(_1031_),
    .C1(_0584_),
    .X(_1032_));
 sky130_fd_sc_hd__mux4_1 _2240_ (.A0(\ram[44][7] ),
    .A1(\ram[45][7] ),
    .A2(\ram[46][7] ),
    .A3(\ram[47][7] ),
    .S0(_0567_),
    .S1(_0728_),
    .X(_1033_));
 sky130_fd_sc_hd__and2_1 _2241_ (.A(_0545_),
    .B(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__and2b_1 _2242_ (.A_N(_0651_),
    .B(\ram[40][7] ),
    .X(_1035_));
 sky130_fd_sc_hd__a21o_1 _2243_ (.A1(_0600_),
    .A2(\ram[41][7] ),
    .B1(_0577_),
    .X(_1036_));
 sky130_fd_sc_hd__mux2_1 _2244_ (.A0(\ram[42][7] ),
    .A1(\ram[43][7] ),
    .S(_0733_),
    .X(_1037_));
 sky130_fd_sc_hd__o221a_1 _2245_ (.A1(_1035_),
    .A2(_1036_),
    .B1(_1037_),
    .B2(_0934_),
    .C1(_0944_),
    .X(_1038_));
 sky130_fd_sc_hd__o21a_1 _2246_ (.A1(_1034_),
    .A2(_1038_),
    .B1(_0542_),
    .X(_1039_));
 sky130_fd_sc_hd__and2b_1 _2247_ (.A_N(_0561_),
    .B(\ram[36][7] ),
    .X(_1040_));
 sky130_fd_sc_hd__a21o_1 _2248_ (.A1(_0568_),
    .A2(\ram[37][7] ),
    .B1(_0577_),
    .X(_1041_));
 sky130_fd_sc_hd__mux2_1 _2249_ (.A0(\ram[38][7] ),
    .A1(\ram[39][7] ),
    .S(_0733_),
    .X(_1042_));
 sky130_fd_sc_hd__o221a_1 _2250_ (.A1(_1040_),
    .A2(_1041_),
    .B1(_1042_),
    .B2(_0934_),
    .C1(_0585_),
    .X(_1043_));
 sky130_fd_sc_hd__mux4_1 _2251_ (.A0(\ram[32][7] ),
    .A1(\ram[33][7] ),
    .A2(\ram[34][7] ),
    .A3(\ram[35][7] ),
    .S0(_0629_),
    .S1(_0550_),
    .X(_1044_));
 sky130_fd_sc_hd__and2_1 _2252_ (.A(_0944_),
    .B(_1044_),
    .X(_1045_));
 sky130_fd_sc_hd__o21ba_1 _2253_ (.A1(_1043_),
    .A2(_1045_),
    .B1_N(_0003_),
    .X(_1046_));
 sky130_fd_sc_hd__o31a_1 _2254_ (.A1(_0581_),
    .A2(_1039_),
    .A3(_1046_),
    .B1(_0005_),
    .X(_1047_));
 sky130_fd_sc_hd__a32o_1 _2255_ (.A1(_0659_),
    .A2(_1004_),
    .A3(_1018_),
    .B1(_1032_),
    .B2(_1047_),
    .X(net23));
 sky130_fd_sc_hd__buf_4 _2256_ (.A(net7),
    .X(_1048_));
 sky130_fd_sc_hd__and3_2 _2257_ (.A(_0530_),
    .B(_0533_),
    .C(_0535_),
    .X(_1049_));
 sky130_fd_sc_hd__inv_2 _2258_ (.A(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__inv_4 _2259_ (.A(net15),
    .Y(_1051_));
 sky130_fd_sc_hd__or4_1 _2260_ (.A(_1051_),
    .B(_0537_),
    .C(net5),
    .D(net6),
    .X(_1052_));
 sky130_fd_sc_hd__clkbuf_8 _2261_ (.A(_1052_),
    .X(_1053_));
 sky130_fd_sc_hd__nor2_4 _2262_ (.A(_1050_),
    .B(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__mux2_1 _2263_ (.A0(net205),
    .A1(_1048_),
    .S(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__clkbuf_1 _2264_ (.A(_1055_),
    .X(_0012_));
 sky130_fd_sc_hd__buf_4 _2265_ (.A(net8),
    .X(_1056_));
 sky130_fd_sc_hd__mux2_1 _2266_ (.A0(net160),
    .A1(_1056_),
    .S(_1054_),
    .X(_1057_));
 sky130_fd_sc_hd__clkbuf_1 _2267_ (.A(_1057_),
    .X(_0013_));
 sky130_fd_sc_hd__buf_4 _2268_ (.A(net9),
    .X(_1058_));
 sky130_fd_sc_hd__mux2_1 _2269_ (.A0(net363),
    .A1(_1058_),
    .S(_1054_),
    .X(_1059_));
 sky130_fd_sc_hd__clkbuf_1 _2270_ (.A(_1059_),
    .X(_0014_));
 sky130_fd_sc_hd__buf_4 _2271_ (.A(net10),
    .X(_1060_));
 sky130_fd_sc_hd__mux2_1 _2272_ (.A0(net289),
    .A1(_1060_),
    .S(_1054_),
    .X(_1061_));
 sky130_fd_sc_hd__clkbuf_1 _2273_ (.A(_1061_),
    .X(_0015_));
 sky130_fd_sc_hd__buf_4 _2274_ (.A(net11),
    .X(_1062_));
 sky130_fd_sc_hd__mux2_1 _2275_ (.A0(net331),
    .A1(_1062_),
    .S(_1054_),
    .X(_1063_));
 sky130_fd_sc_hd__clkbuf_1 _2276_ (.A(_1063_),
    .X(_0016_));
 sky130_fd_sc_hd__clkbuf_4 _2277_ (.A(net12),
    .X(_1064_));
 sky130_fd_sc_hd__mux2_1 _2278_ (.A0(net253),
    .A1(_1064_),
    .S(_1054_),
    .X(_1065_));
 sky130_fd_sc_hd__clkbuf_1 _2279_ (.A(_1065_),
    .X(_0017_));
 sky130_fd_sc_hd__clkbuf_4 _2280_ (.A(net13),
    .X(_1066_));
 sky130_fd_sc_hd__mux2_1 _2281_ (.A0(net327),
    .A1(_1066_),
    .S(_1054_),
    .X(_1067_));
 sky130_fd_sc_hd__clkbuf_1 _2282_ (.A(_1067_),
    .X(_0018_));
 sky130_fd_sc_hd__clkbuf_4 _2283_ (.A(net14),
    .X(_1068_));
 sky130_fd_sc_hd__mux2_1 _2284_ (.A0(net312),
    .A1(_1068_),
    .S(_1054_),
    .X(_1069_));
 sky130_fd_sc_hd__clkbuf_1 _2285_ (.A(_1069_),
    .X(_0019_));
 sky130_fd_sc_hd__clkbuf_4 _2286_ (.A(net7),
    .X(_1070_));
 sky130_fd_sc_hd__and4b_2 _2287_ (.A_N(_0540_),
    .B(net5),
    .C(_0537_),
    .D(net15),
    .X(_1071_));
 sky130_fd_sc_hd__and3b_1 _2288_ (.A_N(_0533_),
    .B(_0535_),
    .C(net1),
    .X(_1072_));
 sky130_fd_sc_hd__nand2_4 _2289_ (.A(_1071_),
    .B(_1072_),
    .Y(_1073_));
 sky130_fd_sc_hd__mux2_1 _2290_ (.A0(_1070_),
    .A1(net484),
    .S(_1073_),
    .X(_1074_));
 sky130_fd_sc_hd__clkbuf_1 _2291_ (.A(_1074_),
    .X(_0020_));
 sky130_fd_sc_hd__clkbuf_4 _2292_ (.A(net8),
    .X(_1075_));
 sky130_fd_sc_hd__mux2_1 _2293_ (.A0(_1075_),
    .A1(net209),
    .S(_1073_),
    .X(_1076_));
 sky130_fd_sc_hd__clkbuf_1 _2294_ (.A(_1076_),
    .X(_0021_));
 sky130_fd_sc_hd__clkbuf_4 _2295_ (.A(net9),
    .X(_1077_));
 sky130_fd_sc_hd__mux2_1 _2296_ (.A0(_1077_),
    .A1(net134),
    .S(_1073_),
    .X(_1078_));
 sky130_fd_sc_hd__clkbuf_1 _2297_ (.A(_1078_),
    .X(_0022_));
 sky130_fd_sc_hd__clkbuf_4 _2298_ (.A(net10),
    .X(_1079_));
 sky130_fd_sc_hd__mux2_1 _2299_ (.A0(_1079_),
    .A1(net219),
    .S(_1073_),
    .X(_1080_));
 sky130_fd_sc_hd__clkbuf_1 _2300_ (.A(_1080_),
    .X(_0023_));
 sky130_fd_sc_hd__clkbuf_4 _2301_ (.A(net11),
    .X(_1081_));
 sky130_fd_sc_hd__mux2_1 _2302_ (.A0(_1081_),
    .A1(net119),
    .S(_1073_),
    .X(_1082_));
 sky130_fd_sc_hd__clkbuf_1 _2303_ (.A(_1082_),
    .X(_0024_));
 sky130_fd_sc_hd__buf_2 _2304_ (.A(net12),
    .X(_1083_));
 sky130_fd_sc_hd__mux2_1 _2305_ (.A0(_1083_),
    .A1(net407),
    .S(_1073_),
    .X(_1084_));
 sky130_fd_sc_hd__clkbuf_1 _2306_ (.A(_1084_),
    .X(_0025_));
 sky130_fd_sc_hd__buf_2 _2307_ (.A(net13),
    .X(_1085_));
 sky130_fd_sc_hd__mux2_1 _2308_ (.A0(_1085_),
    .A1(net404),
    .S(_1073_),
    .X(_1086_));
 sky130_fd_sc_hd__clkbuf_1 _2309_ (.A(_1086_),
    .X(_0026_));
 sky130_fd_sc_hd__buf_2 _2310_ (.A(net14),
    .X(_1087_));
 sky130_fd_sc_hd__mux2_1 _2311_ (.A0(_1087_),
    .A1(net382),
    .S(_1073_),
    .X(_1088_));
 sky130_fd_sc_hd__clkbuf_1 _2312_ (.A(_1088_),
    .X(_0027_));
 sky130_fd_sc_hd__inv_2 _2313_ (.A(net4),
    .Y(_1089_));
 sky130_fd_sc_hd__or3_1 _2314_ (.A(_1089_),
    .B(net5),
    .C(_0540_),
    .X(_1090_));
 sky130_fd_sc_hd__buf_4 _2315_ (.A(_1090_),
    .X(_1091_));
 sky130_fd_sc_hd__or3_4 _2316_ (.A(net1),
    .B(net2),
    .C(net3),
    .X(_1092_));
 sky130_fd_sc_hd__or2_1 _2317_ (.A(_1051_),
    .B(_1092_),
    .X(_1093_));
 sky130_fd_sc_hd__clkbuf_8 _2318_ (.A(_1093_),
    .X(_1094_));
 sky130_fd_sc_hd__nor2_4 _2319_ (.A(_1091_),
    .B(_1094_),
    .Y(_1095_));
 sky130_fd_sc_hd__mux2_1 _2320_ (.A0(net170),
    .A1(_1048_),
    .S(_1095_),
    .X(_1096_));
 sky130_fd_sc_hd__clkbuf_1 _2321_ (.A(_1096_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _2322_ (.A0(net474),
    .A1(_1056_),
    .S(_1095_),
    .X(_1097_));
 sky130_fd_sc_hd__clkbuf_1 _2323_ (.A(_1097_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _2324_ (.A0(net390),
    .A1(_1058_),
    .S(_1095_),
    .X(_1098_));
 sky130_fd_sc_hd__clkbuf_1 _2325_ (.A(_1098_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _2326_ (.A0(net52),
    .A1(_1060_),
    .S(_1095_),
    .X(_1099_));
 sky130_fd_sc_hd__clkbuf_1 _2327_ (.A(_1099_),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _2328_ (.A0(net236),
    .A1(_1062_),
    .S(_1095_),
    .X(_1100_));
 sky130_fd_sc_hd__clkbuf_1 _2329_ (.A(_1100_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _2330_ (.A0(net51),
    .A1(_1064_),
    .S(_1095_),
    .X(_1101_));
 sky130_fd_sc_hd__clkbuf_1 _2331_ (.A(_1101_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _2332_ (.A0(net348),
    .A1(_1066_),
    .S(_1095_),
    .X(_1102_));
 sky130_fd_sc_hd__clkbuf_1 _2333_ (.A(_1102_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _2334_ (.A0(net322),
    .A1(_1068_),
    .S(_1095_),
    .X(_1103_));
 sky130_fd_sc_hd__clkbuf_1 _2335_ (.A(_1103_),
    .X(_0035_));
 sky130_fd_sc_hd__nor2_4 _2336_ (.A(_1053_),
    .B(_1092_),
    .Y(_1104_));
 sky130_fd_sc_hd__mux2_1 _2337_ (.A0(net137),
    .A1(_1048_),
    .S(_1104_),
    .X(_1105_));
 sky130_fd_sc_hd__clkbuf_1 _2338_ (.A(_1105_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _2339_ (.A0(net177),
    .A1(_1056_),
    .S(_1104_),
    .X(_1106_));
 sky130_fd_sc_hd__clkbuf_1 _2340_ (.A(_1106_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _2341_ (.A0(net146),
    .A1(_1058_),
    .S(_1104_),
    .X(_1107_));
 sky130_fd_sc_hd__clkbuf_1 _2342_ (.A(_1107_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _2343_ (.A0(net65),
    .A1(_1060_),
    .S(_1104_),
    .X(_1108_));
 sky130_fd_sc_hd__clkbuf_1 _2344_ (.A(_1108_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _2345_ (.A0(net263),
    .A1(_1062_),
    .S(_1104_),
    .X(_1109_));
 sky130_fd_sc_hd__clkbuf_1 _2346_ (.A(_1109_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _2347_ (.A0(net275),
    .A1(_1064_),
    .S(_1104_),
    .X(_1110_));
 sky130_fd_sc_hd__clkbuf_1 _2348_ (.A(_1110_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _2349_ (.A0(net488),
    .A1(_1066_),
    .S(_1104_),
    .X(_1111_));
 sky130_fd_sc_hd__clkbuf_1 _2350_ (.A(_1111_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _2351_ (.A0(net237),
    .A1(_1068_),
    .S(_1104_),
    .X(_1112_));
 sky130_fd_sc_hd__clkbuf_1 _2352_ (.A(_1112_),
    .X(_0043_));
 sky130_fd_sc_hd__or3b_4 _2353_ (.A(_0530_),
    .B(_0535_),
    .C_N(_0533_),
    .X(_1113_));
 sky130_fd_sc_hd__or2_4 _2354_ (.A(_1051_),
    .B(_1113_),
    .X(_1114_));
 sky130_fd_sc_hd__nor2_4 _2355_ (.A(_1091_),
    .B(_1114_),
    .Y(_1115_));
 sky130_fd_sc_hd__mux2_1 _2356_ (.A0(net392),
    .A1(_1048_),
    .S(_1115_),
    .X(_1116_));
 sky130_fd_sc_hd__clkbuf_1 _2357_ (.A(_1116_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _2358_ (.A0(net277),
    .A1(_1056_),
    .S(_1115_),
    .X(_1117_));
 sky130_fd_sc_hd__clkbuf_1 _2359_ (.A(_1117_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _2360_ (.A0(net297),
    .A1(_1058_),
    .S(_1115_),
    .X(_1118_));
 sky130_fd_sc_hd__clkbuf_1 _2361_ (.A(_1118_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _2362_ (.A0(net313),
    .A1(_1060_),
    .S(_1115_),
    .X(_1119_));
 sky130_fd_sc_hd__clkbuf_1 _2363_ (.A(_1119_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _2364_ (.A0(net309),
    .A1(_1062_),
    .S(_1115_),
    .X(_1120_));
 sky130_fd_sc_hd__clkbuf_1 _2365_ (.A(_1120_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _2366_ (.A0(net94),
    .A1(_1064_),
    .S(_1115_),
    .X(_1121_));
 sky130_fd_sc_hd__clkbuf_1 _2367_ (.A(_1121_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _2368_ (.A0(net242),
    .A1(_1066_),
    .S(_1115_),
    .X(_1122_));
 sky130_fd_sc_hd__clkbuf_1 _2369_ (.A(_1122_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _2370_ (.A0(net178),
    .A1(_1068_),
    .S(_1115_),
    .X(_1123_));
 sky130_fd_sc_hd__clkbuf_1 _2371_ (.A(_1123_),
    .X(_0051_));
 sky130_fd_sc_hd__inv_2 _2372_ (.A(net5),
    .Y(_1124_));
 sky130_fd_sc_hd__and3b_2 _2373_ (.A_N(_0540_),
    .B(_0537_),
    .C(_1124_),
    .X(_1125_));
 sky130_fd_sc_hd__and4b_1 _2374_ (.A_N(_0535_),
    .B(_0533_),
    .C(net15),
    .D(_0530_),
    .X(_1126_));
 sky130_fd_sc_hd__clkbuf_8 _2375_ (.A(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__nand2_4 _2376_ (.A(_1125_),
    .B(_1127_),
    .Y(_1128_));
 sky130_fd_sc_hd__mux2_1 _2377_ (.A0(_1070_),
    .A1(net522),
    .S(_1128_),
    .X(_1129_));
 sky130_fd_sc_hd__clkbuf_1 _2378_ (.A(_1129_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _2379_ (.A0(_1075_),
    .A1(net473),
    .S(_1128_),
    .X(_1130_));
 sky130_fd_sc_hd__clkbuf_1 _2380_ (.A(_1130_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _2381_ (.A0(_1077_),
    .A1(net528),
    .S(_1128_),
    .X(_1131_));
 sky130_fd_sc_hd__clkbuf_1 _2382_ (.A(_1131_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _2383_ (.A0(_1079_),
    .A1(net490),
    .S(_1128_),
    .X(_1132_));
 sky130_fd_sc_hd__clkbuf_1 _2384_ (.A(_1132_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _2385_ (.A0(_1081_),
    .A1(net530),
    .S(_1128_),
    .X(_1133_));
 sky130_fd_sc_hd__clkbuf_1 _2386_ (.A(_1133_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _2387_ (.A0(_1083_),
    .A1(net303),
    .S(_1128_),
    .X(_1134_));
 sky130_fd_sc_hd__clkbuf_1 _2388_ (.A(_1134_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _2389_ (.A0(_1085_),
    .A1(net435),
    .S(_1128_),
    .X(_1135_));
 sky130_fd_sc_hd__clkbuf_1 _2390_ (.A(_1135_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _2391_ (.A0(_1087_),
    .A1(net206),
    .S(_1128_),
    .X(_1136_));
 sky130_fd_sc_hd__clkbuf_1 _2392_ (.A(_1136_),
    .X(_0059_));
 sky130_fd_sc_hd__or3b_4 _2393_ (.A(_0530_),
    .B(_0533_),
    .C_N(_0535_),
    .X(_1137_));
 sky130_fd_sc_hd__or2_4 _2394_ (.A(_1051_),
    .B(_1137_),
    .X(_1138_));
 sky130_fd_sc_hd__nor2_4 _2395_ (.A(_1091_),
    .B(_1138_),
    .Y(_1139_));
 sky130_fd_sc_hd__mux2_1 _2396_ (.A0(net262),
    .A1(_1048_),
    .S(_1139_),
    .X(_1140_));
 sky130_fd_sc_hd__clkbuf_1 _2397_ (.A(_1140_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _2398_ (.A0(net42),
    .A1(_1056_),
    .S(_1139_),
    .X(_1141_));
 sky130_fd_sc_hd__clkbuf_1 _2399_ (.A(_1141_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _2400_ (.A0(net70),
    .A1(_1058_),
    .S(_1139_),
    .X(_1142_));
 sky130_fd_sc_hd__clkbuf_1 _2401_ (.A(_1142_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _2402_ (.A0(net462),
    .A1(_1060_),
    .S(_1139_),
    .X(_1143_));
 sky130_fd_sc_hd__clkbuf_1 _2403_ (.A(_1143_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _2404_ (.A0(net387),
    .A1(_1062_),
    .S(_1139_),
    .X(_1144_));
 sky130_fd_sc_hd__clkbuf_1 _2405_ (.A(_1144_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _2406_ (.A0(net386),
    .A1(_1064_),
    .S(_1139_),
    .X(_1145_));
 sky130_fd_sc_hd__clkbuf_1 _2407_ (.A(_1145_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _2408_ (.A0(net224),
    .A1(_1066_),
    .S(_1139_),
    .X(_1146_));
 sky130_fd_sc_hd__clkbuf_1 _2409_ (.A(_1146_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _2410_ (.A0(net384),
    .A1(_1068_),
    .S(_1139_),
    .X(_1147_));
 sky130_fd_sc_hd__clkbuf_1 _2411_ (.A(_1147_),
    .X(_0067_));
 sky130_fd_sc_hd__and2_1 _2412_ (.A(net15),
    .B(_1072_),
    .X(_1148_));
 sky130_fd_sc_hd__clkbuf_8 _2413_ (.A(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__nand2_4 _2414_ (.A(_1125_),
    .B(_1149_),
    .Y(_1150_));
 sky130_fd_sc_hd__mux2_1 _2415_ (.A0(_1070_),
    .A1(net241),
    .S(_1150_),
    .X(_1151_));
 sky130_fd_sc_hd__clkbuf_1 _2416_ (.A(_1151_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _2417_ (.A0(_1075_),
    .A1(net54),
    .S(_1150_),
    .X(_1152_));
 sky130_fd_sc_hd__clkbuf_1 _2418_ (.A(_1152_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _2419_ (.A0(_1077_),
    .A1(net40),
    .S(_1150_),
    .X(_1153_));
 sky130_fd_sc_hd__clkbuf_1 _2420_ (.A(_1153_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _2421_ (.A0(_1079_),
    .A1(net457),
    .S(_1150_),
    .X(_1154_));
 sky130_fd_sc_hd__clkbuf_1 _2422_ (.A(_1154_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _2423_ (.A0(_1081_),
    .A1(net288),
    .S(_1150_),
    .X(_1155_));
 sky130_fd_sc_hd__clkbuf_1 _2424_ (.A(_1155_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _2425_ (.A0(_1083_),
    .A1(net375),
    .S(_1150_),
    .X(_1156_));
 sky130_fd_sc_hd__clkbuf_1 _2426_ (.A(_1156_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _2427_ (.A0(_1085_),
    .A1(net343),
    .S(_1150_),
    .X(_1157_));
 sky130_fd_sc_hd__clkbuf_1 _2428_ (.A(_1157_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _2429_ (.A0(_1087_),
    .A1(net251),
    .S(_1150_),
    .X(_1158_));
 sky130_fd_sc_hd__clkbuf_1 _2430_ (.A(_1158_),
    .X(_0075_));
 sky130_fd_sc_hd__and3b_1 _2431_ (.A_N(_0530_),
    .B(net2),
    .C(net3),
    .X(_1159_));
 sky130_fd_sc_hd__and2_1 _2432_ (.A(net15),
    .B(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__clkbuf_8 _2433_ (.A(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__nand2_4 _2434_ (.A(_1125_),
    .B(_1161_),
    .Y(_1162_));
 sky130_fd_sc_hd__mux2_1 _2435_ (.A0(_1070_),
    .A1(net419),
    .S(_1162_),
    .X(_1163_));
 sky130_fd_sc_hd__clkbuf_1 _2436_ (.A(_1163_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _2437_ (.A0(_1075_),
    .A1(net212),
    .S(_1162_),
    .X(_1164_));
 sky130_fd_sc_hd__clkbuf_1 _2438_ (.A(_1164_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _2439_ (.A0(_1077_),
    .A1(net109),
    .S(_1162_),
    .X(_1165_));
 sky130_fd_sc_hd__clkbuf_1 _2440_ (.A(_1165_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _2441_ (.A0(_1079_),
    .A1(net430),
    .S(_1162_),
    .X(_1166_));
 sky130_fd_sc_hd__clkbuf_1 _2442_ (.A(_1166_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _2443_ (.A0(_1081_),
    .A1(net230),
    .S(_1162_),
    .X(_1167_));
 sky130_fd_sc_hd__clkbuf_1 _2444_ (.A(_1167_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _2445_ (.A0(_1083_),
    .A1(net437),
    .S(_1162_),
    .X(_1168_));
 sky130_fd_sc_hd__clkbuf_1 _2446_ (.A(_1168_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _2447_ (.A0(_1085_),
    .A1(net161),
    .S(_1162_),
    .X(_1169_));
 sky130_fd_sc_hd__clkbuf_1 _2448_ (.A(_1169_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _2449_ (.A0(_1087_),
    .A1(net421),
    .S(_1162_),
    .X(_1170_));
 sky130_fd_sc_hd__clkbuf_1 _2450_ (.A(_1170_),
    .X(_0083_));
 sky130_fd_sc_hd__nand2_4 _2451_ (.A(net15),
    .B(_1049_),
    .Y(_1171_));
 sky130_fd_sc_hd__nor2_4 _2452_ (.A(_1091_),
    .B(_1171_),
    .Y(_1172_));
 sky130_fd_sc_hd__mux2_1 _2453_ (.A0(net238),
    .A1(_1048_),
    .S(_1172_),
    .X(_1173_));
 sky130_fd_sc_hd__clkbuf_1 _2454_ (.A(_1173_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _2455_ (.A0(net37),
    .A1(_1056_),
    .S(_1172_),
    .X(_1174_));
 sky130_fd_sc_hd__clkbuf_1 _2456_ (.A(_1174_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _2457_ (.A0(net60),
    .A1(_1058_),
    .S(_1172_),
    .X(_1175_));
 sky130_fd_sc_hd__clkbuf_1 _2458_ (.A(_1175_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _2459_ (.A0(net380),
    .A1(_1060_),
    .S(_1172_),
    .X(_1176_));
 sky130_fd_sc_hd__clkbuf_1 _2460_ (.A(_1176_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _2461_ (.A0(net129),
    .A1(_1062_),
    .S(_1172_),
    .X(_1177_));
 sky130_fd_sc_hd__clkbuf_1 _2462_ (.A(_1177_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _2463_ (.A0(net319),
    .A1(_1064_),
    .S(_1172_),
    .X(_1178_));
 sky130_fd_sc_hd__clkbuf_1 _2464_ (.A(_1178_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _2465_ (.A0(net31),
    .A1(_1066_),
    .S(_1172_),
    .X(_1179_));
 sky130_fd_sc_hd__clkbuf_1 _2466_ (.A(_1179_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _2467_ (.A0(net221),
    .A1(_1068_),
    .S(_1172_),
    .X(_1180_));
 sky130_fd_sc_hd__clkbuf_1 _2468_ (.A(_1180_),
    .X(_0091_));
 sky130_fd_sc_hd__clkbuf_4 _2469_ (.A(net7),
    .X(_1181_));
 sky130_fd_sc_hd__or3_1 _2470_ (.A(_0537_),
    .B(_1124_),
    .C(_0540_),
    .X(_1182_));
 sky130_fd_sc_hd__buf_4 _2471_ (.A(_1182_),
    .X(_1183_));
 sky130_fd_sc_hd__nor2_4 _2472_ (.A(_1094_),
    .B(_1183_),
    .Y(_1184_));
 sky130_fd_sc_hd__mux2_1 _2473_ (.A0(net203),
    .A1(_1181_),
    .S(_1184_),
    .X(_1185_));
 sky130_fd_sc_hd__clkbuf_1 _2474_ (.A(_1185_),
    .X(_0092_));
 sky130_fd_sc_hd__buf_2 _2475_ (.A(net8),
    .X(_1186_));
 sky130_fd_sc_hd__mux2_1 _2476_ (.A0(net276),
    .A1(_1186_),
    .S(_1184_),
    .X(_1187_));
 sky130_fd_sc_hd__clkbuf_1 _2477_ (.A(_1187_),
    .X(_0093_));
 sky130_fd_sc_hd__clkbuf_4 _2478_ (.A(net9),
    .X(_1188_));
 sky130_fd_sc_hd__mux2_1 _2479_ (.A0(net64),
    .A1(_1188_),
    .S(_1184_),
    .X(_1189_));
 sky130_fd_sc_hd__clkbuf_1 _2480_ (.A(_1189_),
    .X(_0094_));
 sky130_fd_sc_hd__clkbuf_4 _2481_ (.A(net10),
    .X(_1190_));
 sky130_fd_sc_hd__mux2_1 _2482_ (.A0(net110),
    .A1(_1190_),
    .S(_1184_),
    .X(_1191_));
 sky130_fd_sc_hd__clkbuf_1 _2483_ (.A(_1191_),
    .X(_0095_));
 sky130_fd_sc_hd__clkbuf_4 _2484_ (.A(net11),
    .X(_1192_));
 sky130_fd_sc_hd__mux2_1 _2485_ (.A0(net217),
    .A1(_1192_),
    .S(_1184_),
    .X(_1193_));
 sky130_fd_sc_hd__clkbuf_1 _2486_ (.A(_1193_),
    .X(_0096_));
 sky130_fd_sc_hd__buf_2 _2487_ (.A(net12),
    .X(_1194_));
 sky130_fd_sc_hd__mux2_1 _2488_ (.A0(net186),
    .A1(_1194_),
    .S(_1184_),
    .X(_1195_));
 sky130_fd_sc_hd__clkbuf_1 _2489_ (.A(_1195_),
    .X(_0097_));
 sky130_fd_sc_hd__buf_2 _2490_ (.A(net13),
    .X(_1196_));
 sky130_fd_sc_hd__mux2_1 _2491_ (.A0(net34),
    .A1(_1196_),
    .S(_1184_),
    .X(_1197_));
 sky130_fd_sc_hd__clkbuf_1 _2492_ (.A(_1197_),
    .X(_0098_));
 sky130_fd_sc_hd__clkbuf_4 _2493_ (.A(net14),
    .X(_1198_));
 sky130_fd_sc_hd__mux2_1 _2494_ (.A0(net43),
    .A1(_1198_),
    .S(_1184_),
    .X(_1199_));
 sky130_fd_sc_hd__clkbuf_1 _2495_ (.A(_1199_),
    .X(_0099_));
 sky130_fd_sc_hd__or3b_4 _2496_ (.A(_0533_),
    .B(_0535_),
    .C_N(_0530_),
    .X(_1200_));
 sky130_fd_sc_hd__or2_4 _2497_ (.A(_1051_),
    .B(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__nor2_4 _2498_ (.A(_1183_),
    .B(_1201_),
    .Y(_1202_));
 sky130_fd_sc_hd__mux2_1 _2499_ (.A0(net141),
    .A1(_1181_),
    .S(_1202_),
    .X(_1203_));
 sky130_fd_sc_hd__clkbuf_1 _2500_ (.A(_1203_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _2501_ (.A0(net176),
    .A1(_1186_),
    .S(_1202_),
    .X(_1204_));
 sky130_fd_sc_hd__clkbuf_1 _2502_ (.A(_1204_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _2503_ (.A0(net138),
    .A1(_1188_),
    .S(_1202_),
    .X(_1205_));
 sky130_fd_sc_hd__clkbuf_1 _2504_ (.A(_1205_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _2505_ (.A0(net394),
    .A1(_1190_),
    .S(_1202_),
    .X(_1206_));
 sky130_fd_sc_hd__clkbuf_1 _2506_ (.A(_1206_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _2507_ (.A0(net155),
    .A1(_1192_),
    .S(_1202_),
    .X(_1207_));
 sky130_fd_sc_hd__clkbuf_1 _2508_ (.A(_1207_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _2509_ (.A0(net525),
    .A1(_1194_),
    .S(_1202_),
    .X(_1208_));
 sky130_fd_sc_hd__clkbuf_1 _2510_ (.A(_1208_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _2511_ (.A0(net72),
    .A1(_1196_),
    .S(_1202_),
    .X(_1209_));
 sky130_fd_sc_hd__clkbuf_1 _2512_ (.A(_1209_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _2513_ (.A0(net90),
    .A1(_1198_),
    .S(_1202_),
    .X(_1210_));
 sky130_fd_sc_hd__clkbuf_1 _2514_ (.A(_1210_),
    .X(_0107_));
 sky130_fd_sc_hd__nor2_4 _2515_ (.A(_1114_),
    .B(_1183_),
    .Y(_1211_));
 sky130_fd_sc_hd__mux2_1 _2516_ (.A0(net318),
    .A1(_1181_),
    .S(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__clkbuf_1 _2517_ (.A(_1212_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _2518_ (.A0(net410),
    .A1(_1186_),
    .S(_1211_),
    .X(_1213_));
 sky130_fd_sc_hd__clkbuf_1 _2519_ (.A(_1213_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _2520_ (.A0(net336),
    .A1(_1188_),
    .S(_1211_),
    .X(_1214_));
 sky130_fd_sc_hd__clkbuf_1 _2521_ (.A(_1214_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _2522_ (.A0(net489),
    .A1(_1190_),
    .S(_1211_),
    .X(_1215_));
 sky130_fd_sc_hd__clkbuf_1 _2523_ (.A(_1215_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _2524_ (.A0(net373),
    .A1(_1192_),
    .S(_1211_),
    .X(_1216_));
 sky130_fd_sc_hd__clkbuf_1 _2525_ (.A(_1216_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _2526_ (.A0(net425),
    .A1(_1194_),
    .S(_1211_),
    .X(_1217_));
 sky130_fd_sc_hd__clkbuf_1 _2527_ (.A(_1217_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _2528_ (.A0(net96),
    .A1(_1196_),
    .S(_1211_),
    .X(_1218_));
 sky130_fd_sc_hd__clkbuf_1 _2529_ (.A(_1218_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _2530_ (.A0(net41),
    .A1(_1198_),
    .S(_1211_),
    .X(_1219_));
 sky130_fd_sc_hd__clkbuf_1 _2531_ (.A(_1219_),
    .X(_0115_));
 sky130_fd_sc_hd__nor2_4 _2532_ (.A(_1053_),
    .B(_1200_),
    .Y(_1220_));
 sky130_fd_sc_hd__mux2_1 _2533_ (.A0(net29),
    .A1(_1181_),
    .S(_1220_),
    .X(_1221_));
 sky130_fd_sc_hd__clkbuf_1 _2534_ (.A(_1221_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _2535_ (.A0(net222),
    .A1(_1186_),
    .S(_1220_),
    .X(_1222_));
 sky130_fd_sc_hd__clkbuf_1 _2536_ (.A(_1222_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _2537_ (.A0(net136),
    .A1(_1188_),
    .S(_1220_),
    .X(_1223_));
 sky130_fd_sc_hd__clkbuf_1 _2538_ (.A(_1223_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _2539_ (.A0(net293),
    .A1(_1190_),
    .S(_1220_),
    .X(_1224_));
 sky130_fd_sc_hd__clkbuf_1 _2540_ (.A(_1224_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _2541_ (.A0(net148),
    .A1(_1192_),
    .S(_1220_),
    .X(_1225_));
 sky130_fd_sc_hd__clkbuf_1 _2542_ (.A(_1225_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _2543_ (.A0(net82),
    .A1(_1194_),
    .S(_1220_),
    .X(_1226_));
 sky130_fd_sc_hd__clkbuf_1 _2544_ (.A(_1226_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _2545_ (.A0(net158),
    .A1(_1196_),
    .S(_1220_),
    .X(_1227_));
 sky130_fd_sc_hd__clkbuf_1 _2546_ (.A(_1227_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _2547_ (.A0(net370),
    .A1(_1198_),
    .S(_1220_),
    .X(_1228_));
 sky130_fd_sc_hd__clkbuf_1 _2548_ (.A(_1228_),
    .X(_0123_));
 sky130_fd_sc_hd__nor2_4 _2549_ (.A(_1138_),
    .B(_1183_),
    .Y(_1229_));
 sky130_fd_sc_hd__mux2_1 _2550_ (.A0(net88),
    .A1(_1181_),
    .S(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__clkbuf_1 _2551_ (.A(_1230_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _2552_ (.A0(net338),
    .A1(_1186_),
    .S(_1229_),
    .X(_1231_));
 sky130_fd_sc_hd__clkbuf_1 _2553_ (.A(_1231_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _2554_ (.A0(net49),
    .A1(_1188_),
    .S(_1229_),
    .X(_1232_));
 sky130_fd_sc_hd__clkbuf_1 _2555_ (.A(_1232_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _2556_ (.A0(net130),
    .A1(_1190_),
    .S(_1229_),
    .X(_1233_));
 sky130_fd_sc_hd__clkbuf_1 _2557_ (.A(_1233_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _2558_ (.A0(net84),
    .A1(_1192_),
    .S(_1229_),
    .X(_1234_));
 sky130_fd_sc_hd__clkbuf_1 _2559_ (.A(_1234_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _2560_ (.A0(net311),
    .A1(_1194_),
    .S(_1229_),
    .X(_1235_));
 sky130_fd_sc_hd__clkbuf_1 _2561_ (.A(_1235_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _2562_ (.A0(net326),
    .A1(_1196_),
    .S(_1229_),
    .X(_1236_));
 sky130_fd_sc_hd__clkbuf_1 _2563_ (.A(_1236_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _2564_ (.A0(net169),
    .A1(_1198_),
    .S(_1229_),
    .X(_1237_));
 sky130_fd_sc_hd__clkbuf_1 _2565_ (.A(_1237_),
    .X(_0131_));
 sky130_fd_sc_hd__nor3_4 _2566_ (.A(_0537_),
    .B(_1124_),
    .C(_0540_),
    .Y(_1238_));
 sky130_fd_sc_hd__nand2_4 _2567_ (.A(_1149_),
    .B(_1238_),
    .Y(_1239_));
 sky130_fd_sc_hd__mux2_1 _2568_ (.A0(_1070_),
    .A1(net216),
    .S(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__clkbuf_1 _2569_ (.A(_1240_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _2570_ (.A0(_1075_),
    .A1(net464),
    .S(_1239_),
    .X(_1241_));
 sky130_fd_sc_hd__clkbuf_1 _2571_ (.A(_1241_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _2572_ (.A0(_1077_),
    .A1(net305),
    .S(_1239_),
    .X(_1242_));
 sky130_fd_sc_hd__clkbuf_1 _2573_ (.A(_1242_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _2574_ (.A0(_1079_),
    .A1(net106),
    .S(_1239_),
    .X(_1243_));
 sky130_fd_sc_hd__clkbuf_1 _2575_ (.A(_1243_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _2576_ (.A0(_1081_),
    .A1(net199),
    .S(_1239_),
    .X(_1244_));
 sky130_fd_sc_hd__clkbuf_1 _2577_ (.A(_1244_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _2578_ (.A0(_1083_),
    .A1(net351),
    .S(_1239_),
    .X(_1245_));
 sky130_fd_sc_hd__clkbuf_1 _2579_ (.A(_1245_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _2580_ (.A0(_1085_),
    .A1(net115),
    .S(_1239_),
    .X(_1246_));
 sky130_fd_sc_hd__clkbuf_1 _2581_ (.A(_1246_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _2582_ (.A0(_1087_),
    .A1(net101),
    .S(_1239_),
    .X(_1247_));
 sky130_fd_sc_hd__clkbuf_1 _2583_ (.A(_1247_),
    .X(_0139_));
 sky130_fd_sc_hd__nand2_4 _2584_ (.A(_1161_),
    .B(_1238_),
    .Y(_1248_));
 sky130_fd_sc_hd__mux2_1 _2585_ (.A0(_1070_),
    .A1(net121),
    .S(_1248_),
    .X(_1249_));
 sky130_fd_sc_hd__clkbuf_1 _2586_ (.A(_1249_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _2587_ (.A0(_1075_),
    .A1(net259),
    .S(_1248_),
    .X(_1250_));
 sky130_fd_sc_hd__clkbuf_1 _2588_ (.A(_1250_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _2589_ (.A0(_1077_),
    .A1(net123),
    .S(_1248_),
    .X(_1251_));
 sky130_fd_sc_hd__clkbuf_1 _2590_ (.A(_1251_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _2591_ (.A0(_1079_),
    .A1(net211),
    .S(_1248_),
    .X(_1252_));
 sky130_fd_sc_hd__clkbuf_1 _2592_ (.A(_1252_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _2593_ (.A0(_1081_),
    .A1(net165),
    .S(_1248_),
    .X(_1253_));
 sky130_fd_sc_hd__clkbuf_1 _2594_ (.A(_1253_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _2595_ (.A0(_1083_),
    .A1(net248),
    .S(_1248_),
    .X(_1254_));
 sky130_fd_sc_hd__clkbuf_1 _2596_ (.A(_1254_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _2597_ (.A0(_1085_),
    .A1(net329),
    .S(_1248_),
    .X(_1255_));
 sky130_fd_sc_hd__clkbuf_1 _2598_ (.A(_1255_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _2599_ (.A0(_1087_),
    .A1(net127),
    .S(_1248_),
    .X(_1256_));
 sky130_fd_sc_hd__clkbuf_1 _2600_ (.A(_1256_),
    .X(_0147_));
 sky130_fd_sc_hd__nor2_4 _2601_ (.A(_1171_),
    .B(_1183_),
    .Y(_1257_));
 sky130_fd_sc_hd__mux2_1 _2602_ (.A0(net62),
    .A1(_1181_),
    .S(_1257_),
    .X(_1258_));
 sky130_fd_sc_hd__clkbuf_1 _2603_ (.A(_1258_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _2604_ (.A0(net190),
    .A1(_1186_),
    .S(_1257_),
    .X(_1259_));
 sky130_fd_sc_hd__clkbuf_1 _2605_ (.A(_1259_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _2606_ (.A0(net67),
    .A1(_1188_),
    .S(_1257_),
    .X(_1260_));
 sky130_fd_sc_hd__clkbuf_1 _2607_ (.A(_1260_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _2608_ (.A0(net100),
    .A1(_1190_),
    .S(_1257_),
    .X(_1261_));
 sky130_fd_sc_hd__clkbuf_1 _2609_ (.A(_1261_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _2610_ (.A0(net113),
    .A1(_1192_),
    .S(_1257_),
    .X(_1262_));
 sky130_fd_sc_hd__clkbuf_1 _2611_ (.A(_1262_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _2612_ (.A0(net346),
    .A1(_1194_),
    .S(_1257_),
    .X(_1263_));
 sky130_fd_sc_hd__clkbuf_1 _2613_ (.A(_1263_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _2614_ (.A0(net287),
    .A1(_1196_),
    .S(_1257_),
    .X(_1264_));
 sky130_fd_sc_hd__clkbuf_1 _2615_ (.A(_1264_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _2616_ (.A0(net50),
    .A1(_1198_),
    .S(_1257_),
    .X(_1265_));
 sky130_fd_sc_hd__clkbuf_1 _2617_ (.A(_1265_),
    .X(_0155_));
 sky130_fd_sc_hd__or4_4 _2618_ (.A(_1051_),
    .B(_1089_),
    .C(_1124_),
    .D(_0540_),
    .X(_1266_));
 sky130_fd_sc_hd__nor2_4 _2619_ (.A(_1266_),
    .B(_1092_),
    .Y(_1267_));
 sky130_fd_sc_hd__mux2_1 _2620_ (.A0(net145),
    .A1(_1181_),
    .S(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__clkbuf_1 _2621_ (.A(_1268_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _2622_ (.A0(net244),
    .A1(_1186_),
    .S(_1267_),
    .X(_1269_));
 sky130_fd_sc_hd__clkbuf_1 _2623_ (.A(_1269_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _2624_ (.A0(net513),
    .A1(_1188_),
    .S(_1267_),
    .X(_1270_));
 sky130_fd_sc_hd__clkbuf_1 _2625_ (.A(_1270_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _2626_ (.A0(net381),
    .A1(_1190_),
    .S(_1267_),
    .X(_1271_));
 sky130_fd_sc_hd__clkbuf_1 _2627_ (.A(_1271_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _2628_ (.A0(net174),
    .A1(_1192_),
    .S(_1267_),
    .X(_1272_));
 sky130_fd_sc_hd__clkbuf_1 _2629_ (.A(_1272_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _2630_ (.A0(net166),
    .A1(_1194_),
    .S(_1267_),
    .X(_1273_));
 sky130_fd_sc_hd__clkbuf_1 _2631_ (.A(_1273_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _2632_ (.A0(net39),
    .A1(_1196_),
    .S(_1267_),
    .X(_1274_));
 sky130_fd_sc_hd__clkbuf_1 _2633_ (.A(_1274_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _2634_ (.A0(net301),
    .A1(_1198_),
    .S(_1267_),
    .X(_1275_));
 sky130_fd_sc_hd__clkbuf_1 _2635_ (.A(_1275_),
    .X(_0163_));
 sky130_fd_sc_hd__nor2_4 _2636_ (.A(_1266_),
    .B(_1200_),
    .Y(_1276_));
 sky130_fd_sc_hd__mux2_1 _2637_ (.A0(net376),
    .A1(_1181_),
    .S(_1276_),
    .X(_1277_));
 sky130_fd_sc_hd__clkbuf_1 _2638_ (.A(_1277_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _2639_ (.A0(net335),
    .A1(_1186_),
    .S(_1276_),
    .X(_1278_));
 sky130_fd_sc_hd__clkbuf_1 _2640_ (.A(_1278_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _2641_ (.A0(net365),
    .A1(_1188_),
    .S(_1276_),
    .X(_1279_));
 sky130_fd_sc_hd__clkbuf_1 _2642_ (.A(_1279_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _2643_ (.A0(net426),
    .A1(_1190_),
    .S(_1276_),
    .X(_1280_));
 sky130_fd_sc_hd__clkbuf_1 _2644_ (.A(_1280_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _2645_ (.A0(net468),
    .A1(_1192_),
    .S(_1276_),
    .X(_1281_));
 sky130_fd_sc_hd__clkbuf_1 _2646_ (.A(_1281_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _2647_ (.A0(net347),
    .A1(_1194_),
    .S(_1276_),
    .X(_1282_));
 sky130_fd_sc_hd__clkbuf_1 _2648_ (.A(_1282_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _2649_ (.A0(net215),
    .A1(_1196_),
    .S(_1276_),
    .X(_1283_));
 sky130_fd_sc_hd__clkbuf_1 _2650_ (.A(_1283_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _2651_ (.A0(net36),
    .A1(_1198_),
    .S(_1276_),
    .X(_1284_));
 sky130_fd_sc_hd__clkbuf_1 _2652_ (.A(_1284_),
    .X(_0171_));
 sky130_fd_sc_hd__nor2_4 _2653_ (.A(_1266_),
    .B(_1113_),
    .Y(_1285_));
 sky130_fd_sc_hd__mux2_1 _2654_ (.A0(net184),
    .A1(_1181_),
    .S(_1285_),
    .X(_1286_));
 sky130_fd_sc_hd__clkbuf_1 _2655_ (.A(_1286_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _2656_ (.A0(net140),
    .A1(_1186_),
    .S(_1285_),
    .X(_1287_));
 sky130_fd_sc_hd__clkbuf_1 _2657_ (.A(_1287_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _2658_ (.A0(net261),
    .A1(_1188_),
    .S(_1285_),
    .X(_1288_));
 sky130_fd_sc_hd__clkbuf_1 _2659_ (.A(_1288_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _2660_ (.A0(net149),
    .A1(_1190_),
    .S(_1285_),
    .X(_1289_));
 sky130_fd_sc_hd__clkbuf_1 _2661_ (.A(_1289_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _2662_ (.A0(net153),
    .A1(_1192_),
    .S(_1285_),
    .X(_1290_));
 sky130_fd_sc_hd__clkbuf_1 _2663_ (.A(_1290_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _2664_ (.A0(net198),
    .A1(_1194_),
    .S(_1285_),
    .X(_1291_));
 sky130_fd_sc_hd__clkbuf_1 _2665_ (.A(_1291_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _2666_ (.A0(net260),
    .A1(_1196_),
    .S(_1285_),
    .X(_1292_));
 sky130_fd_sc_hd__clkbuf_1 _2667_ (.A(_1292_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _2668_ (.A0(net226),
    .A1(_1198_),
    .S(_1285_),
    .X(_1293_));
 sky130_fd_sc_hd__clkbuf_1 _2669_ (.A(_1293_),
    .X(_0179_));
 sky130_fd_sc_hd__or4bb_4 _2670_ (.A(_0535_),
    .B(_1266_),
    .C_N(_0530_),
    .D_N(_0533_),
    .X(_1294_));
 sky130_fd_sc_hd__mux2_1 _2671_ (.A0(_1070_),
    .A1(net466),
    .S(_1294_),
    .X(_1295_));
 sky130_fd_sc_hd__clkbuf_1 _2672_ (.A(_1295_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _2673_ (.A0(_1075_),
    .A1(net357),
    .S(_1294_),
    .X(_1296_));
 sky130_fd_sc_hd__clkbuf_1 _2674_ (.A(_1296_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _2675_ (.A0(_1077_),
    .A1(net498),
    .S(_1294_),
    .X(_1297_));
 sky130_fd_sc_hd__clkbuf_1 _2676_ (.A(_1297_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _2677_ (.A0(_1079_),
    .A1(net486),
    .S(_1294_),
    .X(_1298_));
 sky130_fd_sc_hd__clkbuf_1 _2678_ (.A(_1298_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _2679_ (.A0(_1081_),
    .A1(net487),
    .S(_1294_),
    .X(_1299_));
 sky130_fd_sc_hd__clkbuf_1 _2680_ (.A(_1299_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _2681_ (.A0(_1083_),
    .A1(net427),
    .S(_1294_),
    .X(_1300_));
 sky130_fd_sc_hd__clkbuf_1 _2682_ (.A(_1300_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _2683_ (.A0(_1085_),
    .A1(net449),
    .S(_1294_),
    .X(_1301_));
 sky130_fd_sc_hd__clkbuf_1 _2684_ (.A(_1301_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _2685_ (.A0(_1087_),
    .A1(net391),
    .S(_1294_),
    .X(_1302_));
 sky130_fd_sc_hd__clkbuf_1 _2686_ (.A(_1302_),
    .X(_0187_));
 sky130_fd_sc_hd__nor2_4 _2687_ (.A(_1266_),
    .B(_1137_),
    .Y(_1303_));
 sky130_fd_sc_hd__mux2_1 _2688_ (.A0(net118),
    .A1(_1181_),
    .S(_1303_),
    .X(_1304_));
 sky130_fd_sc_hd__clkbuf_1 _2689_ (.A(_1304_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _2690_ (.A0(net256),
    .A1(_1186_),
    .S(_1303_),
    .X(_1305_));
 sky130_fd_sc_hd__clkbuf_1 _2691_ (.A(_1305_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _2692_ (.A0(net91),
    .A1(_1188_),
    .S(_1303_),
    .X(_1306_));
 sky130_fd_sc_hd__clkbuf_1 _2693_ (.A(_1306_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _2694_ (.A0(net66),
    .A1(_1190_),
    .S(_1303_),
    .X(_1307_));
 sky130_fd_sc_hd__clkbuf_1 _2695_ (.A(_1307_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _2696_ (.A0(net75),
    .A1(_1192_),
    .S(_1303_),
    .X(_1308_));
 sky130_fd_sc_hd__clkbuf_1 _2697_ (.A(_1308_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _2698_ (.A0(net409),
    .A1(_1194_),
    .S(_1303_),
    .X(_1309_));
 sky130_fd_sc_hd__clkbuf_1 _2699_ (.A(_1309_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _2700_ (.A0(net102),
    .A1(_1196_),
    .S(_1303_),
    .X(_1310_));
 sky130_fd_sc_hd__clkbuf_1 _2701_ (.A(_1310_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _2702_ (.A0(net128),
    .A1(_1198_),
    .S(_1303_),
    .X(_1311_));
 sky130_fd_sc_hd__clkbuf_1 _2703_ (.A(_1311_),
    .X(_0195_));
 sky130_fd_sc_hd__clkbuf_4 _2704_ (.A(net7),
    .X(_1312_));
 sky130_fd_sc_hd__nor2_4 _2705_ (.A(_1053_),
    .B(_1113_),
    .Y(_1313_));
 sky130_fd_sc_hd__mux2_1 _2706_ (.A0(net218),
    .A1(_1312_),
    .S(_1313_),
    .X(_1314_));
 sky130_fd_sc_hd__clkbuf_1 _2707_ (.A(_1314_),
    .X(_0196_));
 sky130_fd_sc_hd__buf_4 _2708_ (.A(net8),
    .X(_1315_));
 sky130_fd_sc_hd__mux2_1 _2709_ (.A0(net120),
    .A1(_1315_),
    .S(_1313_),
    .X(_1316_));
 sky130_fd_sc_hd__clkbuf_1 _2710_ (.A(_1316_),
    .X(_0197_));
 sky130_fd_sc_hd__buf_4 _2711_ (.A(net9),
    .X(_1317_));
 sky130_fd_sc_hd__mux2_1 _2712_ (.A0(net117),
    .A1(_1317_),
    .S(_1313_),
    .X(_1318_));
 sky130_fd_sc_hd__clkbuf_1 _2713_ (.A(_1318_),
    .X(_0198_));
 sky130_fd_sc_hd__buf_4 _2714_ (.A(net10),
    .X(_1319_));
 sky130_fd_sc_hd__mux2_1 _2715_ (.A0(net114),
    .A1(_1319_),
    .S(_1313_),
    .X(_1320_));
 sky130_fd_sc_hd__clkbuf_1 _2716_ (.A(_1320_),
    .X(_0199_));
 sky130_fd_sc_hd__buf_4 _2717_ (.A(net11),
    .X(_1321_));
 sky130_fd_sc_hd__mux2_1 _2718_ (.A0(net353),
    .A1(_1321_),
    .S(_1313_),
    .X(_1322_));
 sky130_fd_sc_hd__clkbuf_1 _2719_ (.A(_1322_),
    .X(_0200_));
 sky130_fd_sc_hd__buf_4 _2720_ (.A(net12),
    .X(_1323_));
 sky130_fd_sc_hd__mux2_1 _2721_ (.A0(net360),
    .A1(_1323_),
    .S(_1313_),
    .X(_1324_));
 sky130_fd_sc_hd__clkbuf_1 _2722_ (.A(_1324_),
    .X(_0201_));
 sky130_fd_sc_hd__clkbuf_4 _2723_ (.A(net13),
    .X(_1325_));
 sky130_fd_sc_hd__mux2_1 _2724_ (.A0(net163),
    .A1(_1325_),
    .S(_1313_),
    .X(_1326_));
 sky130_fd_sc_hd__clkbuf_1 _2725_ (.A(_1326_),
    .X(_0202_));
 sky130_fd_sc_hd__clkbuf_4 _2726_ (.A(net14),
    .X(_1327_));
 sky130_fd_sc_hd__mux2_1 _2727_ (.A0(net378),
    .A1(_1327_),
    .S(_1313_),
    .X(_1328_));
 sky130_fd_sc_hd__clkbuf_1 _2728_ (.A(_1328_),
    .X(_0203_));
 sky130_fd_sc_hd__nand2_4 _2729_ (.A(_1071_),
    .B(_1159_),
    .Y(_1329_));
 sky130_fd_sc_hd__mux2_1 _2730_ (.A0(_1070_),
    .A1(net266),
    .S(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__clkbuf_1 _2731_ (.A(_1330_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _2732_ (.A0(_1075_),
    .A1(net448),
    .S(_1329_),
    .X(_1331_));
 sky130_fd_sc_hd__clkbuf_1 _2733_ (.A(_1331_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _2734_ (.A0(_1077_),
    .A1(net143),
    .S(_1329_),
    .X(_1332_));
 sky130_fd_sc_hd__clkbuf_1 _2735_ (.A(_1332_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _2736_ (.A0(_1079_),
    .A1(net285),
    .S(_1329_),
    .X(_1333_));
 sky130_fd_sc_hd__clkbuf_1 _2737_ (.A(_1333_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _2738_ (.A0(_1081_),
    .A1(net265),
    .S(_1329_),
    .X(_1334_));
 sky130_fd_sc_hd__clkbuf_1 _2739_ (.A(_1334_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _2740_ (.A0(_1083_),
    .A1(net393),
    .S(_1329_),
    .X(_1335_));
 sky130_fd_sc_hd__clkbuf_1 _2741_ (.A(_1335_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _2742_ (.A0(_1085_),
    .A1(net337),
    .S(_1329_),
    .X(_1336_));
 sky130_fd_sc_hd__clkbuf_1 _2743_ (.A(_1336_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _2744_ (.A0(_1087_),
    .A1(net268),
    .S(_1329_),
    .X(_1337_));
 sky130_fd_sc_hd__clkbuf_1 _2745_ (.A(_1337_),
    .X(_0211_));
 sky130_fd_sc_hd__nand2_4 _2746_ (.A(_1049_),
    .B(_1071_),
    .Y(_1338_));
 sky130_fd_sc_hd__mux2_1 _2747_ (.A0(_1070_),
    .A1(net355),
    .S(_1338_),
    .X(_1339_));
 sky130_fd_sc_hd__clkbuf_1 _2748_ (.A(_1339_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _2749_ (.A0(_1075_),
    .A1(net292),
    .S(_1338_),
    .X(_1340_));
 sky130_fd_sc_hd__clkbuf_1 _2750_ (.A(_1340_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _2751_ (.A0(_1077_),
    .A1(net167),
    .S(_1338_),
    .X(_1341_));
 sky130_fd_sc_hd__clkbuf_1 _2752_ (.A(_1341_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _2753_ (.A0(_1079_),
    .A1(net345),
    .S(_1338_),
    .X(_1342_));
 sky130_fd_sc_hd__clkbuf_1 _2754_ (.A(_1342_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _2755_ (.A0(_1081_),
    .A1(net172),
    .S(_1338_),
    .X(_1343_));
 sky130_fd_sc_hd__clkbuf_1 _2756_ (.A(_1343_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _2757_ (.A0(_1083_),
    .A1(net443),
    .S(_1338_),
    .X(_1344_));
 sky130_fd_sc_hd__clkbuf_1 _2758_ (.A(_1344_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _2759_ (.A0(_1085_),
    .A1(net377),
    .S(_1338_),
    .X(_1345_));
 sky130_fd_sc_hd__clkbuf_1 _2760_ (.A(_1345_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _2761_ (.A0(_1087_),
    .A1(net280),
    .S(_1338_),
    .X(_1346_));
 sky130_fd_sc_hd__clkbuf_1 _2762_ (.A(_1346_),
    .X(_0219_));
 sky130_fd_sc_hd__or3b_1 _2763_ (.A(_0537_),
    .B(net5),
    .C_N(_0540_),
    .X(_1347_));
 sky130_fd_sc_hd__buf_4 _2764_ (.A(_1347_),
    .X(_1348_));
 sky130_fd_sc_hd__nor2_4 _2765_ (.A(_1094_),
    .B(_1348_),
    .Y(_1349_));
 sky130_fd_sc_hd__mux2_1 _2766_ (.A0(net179),
    .A1(_1312_),
    .S(_1349_),
    .X(_1350_));
 sky130_fd_sc_hd__clkbuf_1 _2767_ (.A(_1350_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _2768_ (.A0(net249),
    .A1(_1315_),
    .S(_1349_),
    .X(_1351_));
 sky130_fd_sc_hd__clkbuf_1 _2769_ (.A(_1351_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _2770_ (.A0(net495),
    .A1(_1317_),
    .S(_1349_),
    .X(_1352_));
 sky130_fd_sc_hd__clkbuf_1 _2771_ (.A(_1352_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _2772_ (.A0(net295),
    .A1(_1319_),
    .S(_1349_),
    .X(_1353_));
 sky130_fd_sc_hd__clkbuf_1 _2773_ (.A(_1353_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _2774_ (.A0(net97),
    .A1(_1321_),
    .S(_1349_),
    .X(_1354_));
 sky130_fd_sc_hd__clkbuf_1 _2775_ (.A(_1354_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _2776_ (.A0(net126),
    .A1(_1323_),
    .S(_1349_),
    .X(_1355_));
 sky130_fd_sc_hd__clkbuf_1 _2777_ (.A(_1355_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _2778_ (.A0(net162),
    .A1(_1325_),
    .S(_1349_),
    .X(_1356_));
 sky130_fd_sc_hd__clkbuf_1 _2779_ (.A(_1356_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _2780_ (.A0(net434),
    .A1(_1327_),
    .S(_1349_),
    .X(_1357_));
 sky130_fd_sc_hd__clkbuf_1 _2781_ (.A(_1357_),
    .X(_0227_));
 sky130_fd_sc_hd__nor2_4 _2782_ (.A(_1201_),
    .B(_1348_),
    .Y(_1358_));
 sky130_fd_sc_hd__mux2_1 _2783_ (.A0(net274),
    .A1(_1312_),
    .S(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__clkbuf_1 _2784_ (.A(_1359_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _2785_ (.A0(net116),
    .A1(_1315_),
    .S(_1358_),
    .X(_1360_));
 sky130_fd_sc_hd__clkbuf_1 _2786_ (.A(_1360_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _2787_ (.A0(net349),
    .A1(_1317_),
    .S(_1358_),
    .X(_1361_));
 sky130_fd_sc_hd__clkbuf_1 _2788_ (.A(_1361_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _2789_ (.A0(net187),
    .A1(_1319_),
    .S(_1358_),
    .X(_1362_));
 sky130_fd_sc_hd__clkbuf_1 _2790_ (.A(_1362_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _2791_ (.A0(net330),
    .A1(_1321_),
    .S(_1358_),
    .X(_1363_));
 sky130_fd_sc_hd__clkbuf_1 _2792_ (.A(_1363_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _2793_ (.A0(net55),
    .A1(_1323_),
    .S(_1358_),
    .X(_1364_));
 sky130_fd_sc_hd__clkbuf_1 _2794_ (.A(_1364_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _2795_ (.A0(net202),
    .A1(_1325_),
    .S(_1358_),
    .X(_1365_));
 sky130_fd_sc_hd__clkbuf_1 _2796_ (.A(_1365_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _2797_ (.A0(net239),
    .A1(_1327_),
    .S(_1358_),
    .X(_1366_));
 sky130_fd_sc_hd__clkbuf_1 _2798_ (.A(_1366_),
    .X(_0235_));
 sky130_fd_sc_hd__nor2_4 _2799_ (.A(_1114_),
    .B(_1348_),
    .Y(_1367_));
 sky130_fd_sc_hd__mux2_1 _2800_ (.A0(net433),
    .A1(_1312_),
    .S(_1367_),
    .X(_1368_));
 sky130_fd_sc_hd__clkbuf_1 _2801_ (.A(_1368_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _2802_ (.A0(net270),
    .A1(_1315_),
    .S(_1367_),
    .X(_1369_));
 sky130_fd_sc_hd__clkbuf_1 _2803_ (.A(_1369_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _2804_ (.A0(net284),
    .A1(_1317_),
    .S(_1367_),
    .X(_1370_));
 sky130_fd_sc_hd__clkbuf_1 _2805_ (.A(_1370_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _2806_ (.A0(net371),
    .A1(_1319_),
    .S(_1367_),
    .X(_1371_));
 sky130_fd_sc_hd__clkbuf_1 _2807_ (.A(_1371_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _2808_ (.A0(net352),
    .A1(_1321_),
    .S(_1367_),
    .X(_1372_));
 sky130_fd_sc_hd__clkbuf_1 _2809_ (.A(_1372_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _2810_ (.A0(net56),
    .A1(_1323_),
    .S(_1367_),
    .X(_1373_));
 sky130_fd_sc_hd__clkbuf_1 _2811_ (.A(_1373_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _2812_ (.A0(net81),
    .A1(_1325_),
    .S(_1367_),
    .X(_1374_));
 sky130_fd_sc_hd__clkbuf_1 _2813_ (.A(_1374_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _2814_ (.A0(net59),
    .A1(_1327_),
    .S(_1367_),
    .X(_1375_));
 sky130_fd_sc_hd__clkbuf_1 _2815_ (.A(_1375_),
    .X(_0243_));
 sky130_fd_sc_hd__and3_4 _2816_ (.A(_1089_),
    .B(_1124_),
    .C(_0540_),
    .X(_1376_));
 sky130_fd_sc_hd__nand2_4 _2817_ (.A(_1127_),
    .B(_1376_),
    .Y(_1377_));
 sky130_fd_sc_hd__mux2_1 _2818_ (.A0(_1070_),
    .A1(net507),
    .S(_1377_),
    .X(_1378_));
 sky130_fd_sc_hd__clkbuf_1 _2819_ (.A(_1378_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _2820_ (.A0(_1075_),
    .A1(\ram[35][1] ),
    .S(_1377_),
    .X(_1379_));
 sky130_fd_sc_hd__clkbuf_1 _2821_ (.A(_1379_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _2822_ (.A0(_1077_),
    .A1(\ram[35][2] ),
    .S(_1377_),
    .X(_1380_));
 sky130_fd_sc_hd__clkbuf_1 _2823_ (.A(_1380_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _2824_ (.A0(_1079_),
    .A1(net506),
    .S(_1377_),
    .X(_1381_));
 sky130_fd_sc_hd__clkbuf_1 _2825_ (.A(_1381_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _2826_ (.A0(_1081_),
    .A1(net502),
    .S(_1377_),
    .X(_1382_));
 sky130_fd_sc_hd__clkbuf_1 _2827_ (.A(_1382_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _2828_ (.A0(_1083_),
    .A1(net245),
    .S(_1377_),
    .X(_1383_));
 sky130_fd_sc_hd__clkbuf_1 _2829_ (.A(_1383_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _2830_ (.A0(_1085_),
    .A1(net445),
    .S(_1377_),
    .X(_1384_));
 sky130_fd_sc_hd__clkbuf_1 _2831_ (.A(_1384_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _2832_ (.A0(_1087_),
    .A1(net472),
    .S(_1377_),
    .X(_1385_));
 sky130_fd_sc_hd__clkbuf_1 _2833_ (.A(_1385_),
    .X(_0251_));
 sky130_fd_sc_hd__nor2_4 _2834_ (.A(_1138_),
    .B(_1348_),
    .Y(_1386_));
 sky130_fd_sc_hd__mux2_1 _2835_ (.A0(net183),
    .A1(_1312_),
    .S(_1386_),
    .X(_1387_));
 sky130_fd_sc_hd__clkbuf_1 _2836_ (.A(_1387_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _2837_ (.A0(net112),
    .A1(_1315_),
    .S(_1386_),
    .X(_1388_));
 sky130_fd_sc_hd__clkbuf_1 _2838_ (.A(_1388_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _2839_ (.A0(net307),
    .A1(_1317_),
    .S(_1386_),
    .X(_1389_));
 sky130_fd_sc_hd__clkbuf_1 _2840_ (.A(_1389_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _2841_ (.A0(net452),
    .A1(_1319_),
    .S(_1386_),
    .X(_1390_));
 sky130_fd_sc_hd__clkbuf_1 _2842_ (.A(_1390_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _2843_ (.A0(net93),
    .A1(_1321_),
    .S(_1386_),
    .X(_1391_));
 sky130_fd_sc_hd__clkbuf_1 _2844_ (.A(_1391_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _2845_ (.A0(net201),
    .A1(_1323_),
    .S(_1386_),
    .X(_1392_));
 sky130_fd_sc_hd__clkbuf_1 _2846_ (.A(_1392_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _2847_ (.A0(net132),
    .A1(_1325_),
    .S(_1386_),
    .X(_1393_));
 sky130_fd_sc_hd__clkbuf_1 _2848_ (.A(_1393_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _2849_ (.A0(net213),
    .A1(_1327_),
    .S(_1386_),
    .X(_1394_));
 sky130_fd_sc_hd__clkbuf_1 _2850_ (.A(_1394_),
    .X(_0259_));
 sky130_fd_sc_hd__clkbuf_4 _2851_ (.A(net7),
    .X(_1395_));
 sky130_fd_sc_hd__nand2_4 _2852_ (.A(_1149_),
    .B(_1376_),
    .Y(_1396_));
 sky130_fd_sc_hd__mux2_1 _2853_ (.A0(_1395_),
    .A1(\ram[37][0] ),
    .S(_1396_),
    .X(_1397_));
 sky130_fd_sc_hd__clkbuf_1 _2854_ (.A(_1397_),
    .X(_0260_));
 sky130_fd_sc_hd__clkbuf_4 _2855_ (.A(net8),
    .X(_1398_));
 sky130_fd_sc_hd__mux2_1 _2856_ (.A0(_1398_),
    .A1(net517),
    .S(_1396_),
    .X(_1399_));
 sky130_fd_sc_hd__clkbuf_1 _2857_ (.A(_1399_),
    .X(_0261_));
 sky130_fd_sc_hd__clkbuf_4 _2858_ (.A(net9),
    .X(_1400_));
 sky130_fd_sc_hd__mux2_1 _2859_ (.A0(_1400_),
    .A1(net104),
    .S(_1396_),
    .X(_1401_));
 sky130_fd_sc_hd__clkbuf_1 _2860_ (.A(_1401_),
    .X(_0262_));
 sky130_fd_sc_hd__clkbuf_4 _2861_ (.A(net10),
    .X(_1402_));
 sky130_fd_sc_hd__mux2_1 _2862_ (.A0(_1402_),
    .A1(net95),
    .S(_1396_),
    .X(_1403_));
 sky130_fd_sc_hd__clkbuf_1 _2863_ (.A(_1403_),
    .X(_0263_));
 sky130_fd_sc_hd__buf_2 _2864_ (.A(net11),
    .X(_1404_));
 sky130_fd_sc_hd__mux2_1 _2865_ (.A0(_1404_),
    .A1(net477),
    .S(_1396_),
    .X(_1405_));
 sky130_fd_sc_hd__clkbuf_1 _2866_ (.A(_1405_),
    .X(_0264_));
 sky130_fd_sc_hd__buf_2 _2867_ (.A(net12),
    .X(_1406_));
 sky130_fd_sc_hd__mux2_1 _2868_ (.A0(_1406_),
    .A1(net271),
    .S(_1396_),
    .X(_1407_));
 sky130_fd_sc_hd__clkbuf_1 _2869_ (.A(_1407_),
    .X(_0265_));
 sky130_fd_sc_hd__buf_2 _2870_ (.A(net13),
    .X(_1408_));
 sky130_fd_sc_hd__mux2_1 _2871_ (.A0(_1408_),
    .A1(net48),
    .S(_1396_),
    .X(_1409_));
 sky130_fd_sc_hd__clkbuf_1 _2872_ (.A(_1409_),
    .X(_0266_));
 sky130_fd_sc_hd__buf_2 _2873_ (.A(net14),
    .X(_1410_));
 sky130_fd_sc_hd__mux2_1 _2874_ (.A0(_1410_),
    .A1(net500),
    .S(_1396_),
    .X(_1411_));
 sky130_fd_sc_hd__clkbuf_1 _2875_ (.A(_1411_),
    .X(_0267_));
 sky130_fd_sc_hd__nand2_4 _2876_ (.A(_1161_),
    .B(_1376_),
    .Y(_1412_));
 sky130_fd_sc_hd__mux2_1 _2877_ (.A0(_1395_),
    .A1(net316),
    .S(_1412_),
    .X(_1413_));
 sky130_fd_sc_hd__clkbuf_1 _2878_ (.A(_1413_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _2879_ (.A0(_1398_),
    .A1(net453),
    .S(_1412_),
    .X(_1414_));
 sky130_fd_sc_hd__clkbuf_1 _2880_ (.A(_1414_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _2881_ (.A0(_1400_),
    .A1(net142),
    .S(_1412_),
    .X(_1415_));
 sky130_fd_sc_hd__clkbuf_1 _2882_ (.A(_1415_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _2883_ (.A0(_1402_),
    .A1(net58),
    .S(_1412_),
    .X(_1416_));
 sky130_fd_sc_hd__clkbuf_1 _2884_ (.A(_1416_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _2885_ (.A0(_1404_),
    .A1(net291),
    .S(_1412_),
    .X(_1417_));
 sky130_fd_sc_hd__clkbuf_1 _2886_ (.A(_1417_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _2887_ (.A0(_1406_),
    .A1(net369),
    .S(_1412_),
    .X(_1418_));
 sky130_fd_sc_hd__clkbuf_1 _2888_ (.A(_1418_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _2889_ (.A0(_1408_),
    .A1(net45),
    .S(_1412_),
    .X(_1419_));
 sky130_fd_sc_hd__clkbuf_1 _2890_ (.A(_1419_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _2891_ (.A0(_1410_),
    .A1(net389),
    .S(_1412_),
    .X(_1420_));
 sky130_fd_sc_hd__clkbuf_1 _2892_ (.A(_1420_),
    .X(_0275_));
 sky130_fd_sc_hd__and4bb_4 _2893_ (.A_N(_0535_),
    .B_N(_1053_),
    .C(_0530_),
    .D(_0533_),
    .X(_1421_));
 sky130_fd_sc_hd__mux2_1 _2894_ (.A0(net77),
    .A1(_1312_),
    .S(_1421_),
    .X(_1422_));
 sky130_fd_sc_hd__clkbuf_1 _2895_ (.A(_1422_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _2896_ (.A0(net412),
    .A1(_1315_),
    .S(_1421_),
    .X(_1423_));
 sky130_fd_sc_hd__clkbuf_1 _2897_ (.A(_1423_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _2898_ (.A0(net135),
    .A1(_1317_),
    .S(_1421_),
    .X(_1424_));
 sky130_fd_sc_hd__clkbuf_1 _2899_ (.A(_1424_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _2900_ (.A0(net214),
    .A1(_1319_),
    .S(_1421_),
    .X(_1425_));
 sky130_fd_sc_hd__clkbuf_1 _2901_ (.A(_1425_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _2902_ (.A0(net257),
    .A1(_1321_),
    .S(_1421_),
    .X(_1426_));
 sky130_fd_sc_hd__clkbuf_1 _2903_ (.A(_1426_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _2904_ (.A0(net192),
    .A1(_1323_),
    .S(_1421_),
    .X(_1427_));
 sky130_fd_sc_hd__clkbuf_1 _2905_ (.A(_1427_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _2906_ (.A0(net164),
    .A1(_1325_),
    .S(_1421_),
    .X(_1428_));
 sky130_fd_sc_hd__clkbuf_1 _2907_ (.A(_1428_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _2908_ (.A0(net220),
    .A1(_1327_),
    .S(_1421_),
    .X(_1429_));
 sky130_fd_sc_hd__clkbuf_1 _2909_ (.A(_1429_),
    .X(_0283_));
 sky130_fd_sc_hd__and3b_1 _2910_ (.A_N(net5),
    .B(net6),
    .C(_0537_),
    .X(_1430_));
 sky130_fd_sc_hd__buf_6 _2911_ (.A(_1430_),
    .X(_1431_));
 sky130_fd_sc_hd__nor2b_4 _2912_ (.A(_1094_),
    .B_N(_1431_),
    .Y(_1432_));
 sky130_fd_sc_hd__mux2_1 _2913_ (.A0(net125),
    .A1(_1312_),
    .S(_1432_),
    .X(_1433_));
 sky130_fd_sc_hd__clkbuf_1 _2914_ (.A(_1433_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _2915_ (.A0(net328),
    .A1(_1315_),
    .S(_1432_),
    .X(_1434_));
 sky130_fd_sc_hd__clkbuf_1 _2916_ (.A(_1434_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _2917_ (.A0(net299),
    .A1(_1317_),
    .S(_1432_),
    .X(_1435_));
 sky130_fd_sc_hd__clkbuf_1 _2918_ (.A(_1435_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _2919_ (.A0(net196),
    .A1(_1319_),
    .S(_1432_),
    .X(_1436_));
 sky130_fd_sc_hd__clkbuf_1 _2920_ (.A(_1436_),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _2921_ (.A0(net308),
    .A1(_1321_),
    .S(_1432_),
    .X(_1437_));
 sky130_fd_sc_hd__clkbuf_1 _2922_ (.A(_1437_),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _2923_ (.A0(net207),
    .A1(_1323_),
    .S(_1432_),
    .X(_1438_));
 sky130_fd_sc_hd__clkbuf_1 _2924_ (.A(_1438_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _2925_ (.A0(net25),
    .A1(_1325_),
    .S(_1432_),
    .X(_1439_));
 sky130_fd_sc_hd__clkbuf_1 _2926_ (.A(_1439_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _2927_ (.A0(net152),
    .A1(_1327_),
    .S(_1432_),
    .X(_1440_));
 sky130_fd_sc_hd__clkbuf_1 _2928_ (.A(_1440_),
    .X(_0291_));
 sky130_fd_sc_hd__nor2_4 _2929_ (.A(_1051_),
    .B(_1200_),
    .Y(_1441_));
 sky130_fd_sc_hd__nand2_4 _2930_ (.A(_1441_),
    .B(_1431_),
    .Y(_1442_));
 sky130_fd_sc_hd__mux2_1 _2931_ (.A0(_1395_),
    .A1(net47),
    .S(_1442_),
    .X(_1443_));
 sky130_fd_sc_hd__clkbuf_1 _2932_ (.A(_1443_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _2933_ (.A0(_1398_),
    .A1(net340),
    .S(_1442_),
    .X(_1444_));
 sky130_fd_sc_hd__clkbuf_1 _2934_ (.A(_1444_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _2935_ (.A0(_1400_),
    .A1(net304),
    .S(_1442_),
    .X(_1445_));
 sky130_fd_sc_hd__clkbuf_1 _2936_ (.A(_1445_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _2937_ (.A0(_1402_),
    .A1(net26),
    .S(_1442_),
    .X(_1446_));
 sky130_fd_sc_hd__clkbuf_1 _2938_ (.A(_1446_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _2939_ (.A0(_1404_),
    .A1(net83),
    .S(_1442_),
    .X(_1447_));
 sky130_fd_sc_hd__clkbuf_1 _2940_ (.A(_1447_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _2941_ (.A0(_1406_),
    .A1(net27),
    .S(_1442_),
    .X(_1448_));
 sky130_fd_sc_hd__clkbuf_1 _2942_ (.A(_1448_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _2943_ (.A0(_1408_),
    .A1(net99),
    .S(_1442_),
    .X(_1449_));
 sky130_fd_sc_hd__clkbuf_1 _2944_ (.A(_1449_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _2945_ (.A0(_1410_),
    .A1(net32),
    .S(_1442_),
    .X(_1450_));
 sky130_fd_sc_hd__clkbuf_1 _2946_ (.A(_1450_),
    .X(_0299_));
 sky130_fd_sc_hd__nor2_4 _2947_ (.A(_1051_),
    .B(_1113_),
    .Y(_1451_));
 sky130_fd_sc_hd__nand2_4 _2948_ (.A(_1451_),
    .B(_1431_),
    .Y(_1452_));
 sky130_fd_sc_hd__mux2_1 _2949_ (.A0(_1395_),
    .A1(net354),
    .S(_1452_),
    .X(_1453_));
 sky130_fd_sc_hd__clkbuf_1 _2950_ (.A(_1453_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _2951_ (.A0(_1398_),
    .A1(net395),
    .S(_1452_),
    .X(_1454_));
 sky130_fd_sc_hd__clkbuf_1 _2952_ (.A(_1454_),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _2953_ (.A0(_1400_),
    .A1(net273),
    .S(_1452_),
    .X(_1455_));
 sky130_fd_sc_hd__clkbuf_1 _2954_ (.A(_1455_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _2955_ (.A0(_1402_),
    .A1(net456),
    .S(_1452_),
    .X(_1456_));
 sky130_fd_sc_hd__clkbuf_1 _2956_ (.A(_1456_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _2957_ (.A0(_1404_),
    .A1(net469),
    .S(_1452_),
    .X(_1457_));
 sky130_fd_sc_hd__clkbuf_1 _2958_ (.A(_1457_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _2959_ (.A0(_1406_),
    .A1(net200),
    .S(_1452_),
    .X(_1458_));
 sky130_fd_sc_hd__clkbuf_1 _2960_ (.A(_1458_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _2961_ (.A0(_1408_),
    .A1(net333),
    .S(_1452_),
    .X(_1459_));
 sky130_fd_sc_hd__clkbuf_1 _2962_ (.A(_1459_),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _2963_ (.A0(_1410_),
    .A1(net78),
    .S(_1452_),
    .X(_1460_));
 sky130_fd_sc_hd__clkbuf_1 _2964_ (.A(_1460_),
    .X(_0307_));
 sky130_fd_sc_hd__nand2_4 _2965_ (.A(_1127_),
    .B(_1431_),
    .Y(_1461_));
 sky130_fd_sc_hd__mux2_1 _2966_ (.A0(_1395_),
    .A1(net520),
    .S(_1461_),
    .X(_1462_));
 sky130_fd_sc_hd__clkbuf_1 _2967_ (.A(_1462_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _2968_ (.A0(_1398_),
    .A1(net440),
    .S(_1461_),
    .X(_1463_));
 sky130_fd_sc_hd__clkbuf_1 _2969_ (.A(_1463_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _2970_ (.A0(_1400_),
    .A1(net446),
    .S(_1461_),
    .X(_1464_));
 sky130_fd_sc_hd__clkbuf_1 _2971_ (.A(_1464_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _2972_ (.A0(_1402_),
    .A1(net359),
    .S(_1461_),
    .X(_1465_));
 sky130_fd_sc_hd__clkbuf_1 _2973_ (.A(_1465_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _2974_ (.A0(_1404_),
    .A1(net508),
    .S(_1461_),
    .X(_1466_));
 sky130_fd_sc_hd__clkbuf_1 _2975_ (.A(_1466_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _2976_ (.A0(_1406_),
    .A1(net324),
    .S(_1461_),
    .X(_1467_));
 sky130_fd_sc_hd__clkbuf_1 _2977_ (.A(_1467_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _2978_ (.A0(_1408_),
    .A1(net252),
    .S(_1461_),
    .X(_1468_));
 sky130_fd_sc_hd__clkbuf_1 _2979_ (.A(_1468_),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _2980_ (.A0(_1410_),
    .A1(net189),
    .S(_1461_),
    .X(_1469_));
 sky130_fd_sc_hd__clkbuf_1 _2981_ (.A(_1469_),
    .X(_0315_));
 sky130_fd_sc_hd__nor2_4 _2982_ (.A(_1051_),
    .B(_1137_),
    .Y(_1470_));
 sky130_fd_sc_hd__nand2_4 _2983_ (.A(_1470_),
    .B(_1431_),
    .Y(_1471_));
 sky130_fd_sc_hd__mux2_1 _2984_ (.A0(_1395_),
    .A1(net475),
    .S(_1471_),
    .X(_1472_));
 sky130_fd_sc_hd__clkbuf_1 _2985_ (.A(_1472_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _2986_ (.A0(_1398_),
    .A1(net471),
    .S(_1471_),
    .X(_1473_));
 sky130_fd_sc_hd__clkbuf_1 _2987_ (.A(_1473_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _2988_ (.A0(_1400_),
    .A1(net523),
    .S(_1471_),
    .X(_1474_));
 sky130_fd_sc_hd__clkbuf_1 _2989_ (.A(_1474_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _2990_ (.A0(_1402_),
    .A1(net482),
    .S(_1471_),
    .X(_1475_));
 sky130_fd_sc_hd__clkbuf_1 _2991_ (.A(_1475_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _2992_ (.A0(_1404_),
    .A1(net519),
    .S(_1471_),
    .X(_1476_));
 sky130_fd_sc_hd__clkbuf_1 _2993_ (.A(_1476_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _2994_ (.A0(_1406_),
    .A1(net92),
    .S(_1471_),
    .X(_1477_));
 sky130_fd_sc_hd__clkbuf_1 _2995_ (.A(_1477_),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _2996_ (.A0(_1408_),
    .A1(net157),
    .S(_1471_),
    .X(_1478_));
 sky130_fd_sc_hd__clkbuf_1 _2997_ (.A(_1478_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _2998_ (.A0(_1410_),
    .A1(net185),
    .S(_1471_),
    .X(_1479_));
 sky130_fd_sc_hd__clkbuf_1 _2999_ (.A(_1479_),
    .X(_0323_));
 sky130_fd_sc_hd__nand2_4 _3000_ (.A(_1149_),
    .B(_1431_),
    .Y(_1480_));
 sky130_fd_sc_hd__mux2_1 _3001_ (.A0(_1395_),
    .A1(net518),
    .S(_1480_),
    .X(_1481_));
 sky130_fd_sc_hd__clkbuf_1 _3002_ (.A(_1481_),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _3003_ (.A0(_1398_),
    .A1(net470),
    .S(_1480_),
    .X(_1482_));
 sky130_fd_sc_hd__clkbuf_1 _3004_ (.A(_1482_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _3005_ (.A0(_1400_),
    .A1(net501),
    .S(_1480_),
    .X(_1483_));
 sky130_fd_sc_hd__clkbuf_1 _3006_ (.A(_1483_),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _3007_ (.A0(_1402_),
    .A1(net481),
    .S(_1480_),
    .X(_1484_));
 sky130_fd_sc_hd__clkbuf_1 _3008_ (.A(_1484_),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _3009_ (.A0(_1404_),
    .A1(net428),
    .S(_1480_),
    .X(_1485_));
 sky130_fd_sc_hd__clkbuf_1 _3010_ (.A(_1485_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _3011_ (.A0(_1406_),
    .A1(net63),
    .S(_1480_),
    .X(_1486_));
 sky130_fd_sc_hd__clkbuf_1 _3012_ (.A(_1486_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _3013_ (.A0(_1408_),
    .A1(net512),
    .S(_1480_),
    .X(_1487_));
 sky130_fd_sc_hd__clkbuf_1 _3014_ (.A(_1487_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _3015_ (.A0(_1410_),
    .A1(net368),
    .S(_1480_),
    .X(_1488_));
 sky130_fd_sc_hd__clkbuf_1 _3016_ (.A(_1488_),
    .X(_0331_));
 sky130_fd_sc_hd__nand2_4 _3017_ (.A(_1161_),
    .B(_1431_),
    .Y(_1489_));
 sky130_fd_sc_hd__mux2_1 _3018_ (.A0(_1395_),
    .A1(net505),
    .S(_1489_),
    .X(_1490_));
 sky130_fd_sc_hd__clkbuf_1 _3019_ (.A(_1490_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _3020_ (.A0(_1398_),
    .A1(net383),
    .S(_1489_),
    .X(_1491_));
 sky130_fd_sc_hd__clkbuf_1 _3021_ (.A(_1491_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _3022_ (.A0(_1400_),
    .A1(net444),
    .S(_1489_),
    .X(_1492_));
 sky130_fd_sc_hd__clkbuf_1 _3023_ (.A(_1492_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _3024_ (.A0(_1402_),
    .A1(net514),
    .S(_1489_),
    .X(_1493_));
 sky130_fd_sc_hd__clkbuf_1 _3025_ (.A(_1493_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _3026_ (.A0(_1404_),
    .A1(net485),
    .S(_1489_),
    .X(_1494_));
 sky130_fd_sc_hd__clkbuf_1 _3027_ (.A(_1494_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _3028_ (.A0(_1406_),
    .A1(net139),
    .S(_1489_),
    .X(_1495_));
 sky130_fd_sc_hd__clkbuf_1 _3029_ (.A(_1495_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _3030_ (.A0(_1408_),
    .A1(net402),
    .S(_1489_),
    .X(_1496_));
 sky130_fd_sc_hd__clkbuf_1 _3031_ (.A(_1496_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _3032_ (.A0(_1410_),
    .A1(net320),
    .S(_1489_),
    .X(_1497_));
 sky130_fd_sc_hd__clkbuf_1 _3033_ (.A(_1497_),
    .X(_0339_));
 sky130_fd_sc_hd__nor2_4 _3034_ (.A(_1051_),
    .B(_1050_),
    .Y(_1498_));
 sky130_fd_sc_hd__nand2_4 _3035_ (.A(_1498_),
    .B(_1431_),
    .Y(_1499_));
 sky130_fd_sc_hd__mux2_1 _3036_ (.A0(_1395_),
    .A1(net516),
    .S(_1499_),
    .X(_1500_));
 sky130_fd_sc_hd__clkbuf_1 _3037_ (.A(_1500_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _3038_ (.A0(_1398_),
    .A1(net321),
    .S(_1499_),
    .X(_1501_));
 sky130_fd_sc_hd__clkbuf_1 _3039_ (.A(_1501_),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _3040_ (.A0(_1400_),
    .A1(net510),
    .S(_1499_),
    .X(_1502_));
 sky130_fd_sc_hd__clkbuf_1 _3041_ (.A(_1502_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _3042_ (.A0(_1402_),
    .A1(net526),
    .S(_1499_),
    .X(_1503_));
 sky130_fd_sc_hd__clkbuf_1 _3043_ (.A(_1503_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _3044_ (.A0(_1404_),
    .A1(net509),
    .S(_1499_),
    .X(_1504_));
 sky130_fd_sc_hd__clkbuf_1 _3045_ (.A(_1504_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _3046_ (.A0(_1406_),
    .A1(net180),
    .S(_1499_),
    .X(_1505_));
 sky130_fd_sc_hd__clkbuf_1 _3047_ (.A(_1505_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _3048_ (.A0(_1408_),
    .A1(net122),
    .S(_1499_),
    .X(_1506_));
 sky130_fd_sc_hd__clkbuf_1 _3049_ (.A(_1506_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _3050_ (.A0(_1410_),
    .A1(net247),
    .S(_1499_),
    .X(_1507_));
 sky130_fd_sc_hd__clkbuf_1 _3051_ (.A(_1507_),
    .X(_0347_));
 sky130_fd_sc_hd__and3_1 _3052_ (.A(_1089_),
    .B(net5),
    .C(net6),
    .X(_1508_));
 sky130_fd_sc_hd__buf_6 _3053_ (.A(_1508_),
    .X(_1509_));
 sky130_fd_sc_hd__nor2b_4 _3054_ (.A(_1094_),
    .B_N(_1509_),
    .Y(_1510_));
 sky130_fd_sc_hd__mux2_1 _3055_ (.A0(net406),
    .A1(_1312_),
    .S(_1510_),
    .X(_1511_));
 sky130_fd_sc_hd__clkbuf_1 _3056_ (.A(_1511_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _3057_ (.A0(net105),
    .A1(_1315_),
    .S(_1510_),
    .X(_1512_));
 sky130_fd_sc_hd__clkbuf_1 _3058_ (.A(_1512_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _3059_ (.A0(net422),
    .A1(_1317_),
    .S(_1510_),
    .X(_1513_));
 sky130_fd_sc_hd__clkbuf_1 _3060_ (.A(_1513_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _3061_ (.A0(net323),
    .A1(_1319_),
    .S(_1510_),
    .X(_1514_));
 sky130_fd_sc_hd__clkbuf_1 _3062_ (.A(_1514_),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _3063_ (.A0(net272),
    .A1(_1321_),
    .S(_1510_),
    .X(_1515_));
 sky130_fd_sc_hd__clkbuf_1 _3064_ (.A(_1515_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _3065_ (.A0(net87),
    .A1(_1323_),
    .S(_1510_),
    .X(_1516_));
 sky130_fd_sc_hd__clkbuf_1 _3066_ (.A(_1516_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _3067_ (.A0(net61),
    .A1(_1325_),
    .S(_1510_),
    .X(_1517_));
 sky130_fd_sc_hd__clkbuf_1 _3068_ (.A(_1517_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _3069_ (.A0(net38),
    .A1(_1327_),
    .S(_1510_),
    .X(_1518_));
 sky130_fd_sc_hd__clkbuf_1 _3070_ (.A(_1518_),
    .X(_0355_));
 sky130_fd_sc_hd__nor2_4 _3071_ (.A(_1053_),
    .B(_1137_),
    .Y(_1519_));
 sky130_fd_sc_hd__mux2_1 _3072_ (.A0(net258),
    .A1(_1312_),
    .S(_1519_),
    .X(_1520_));
 sky130_fd_sc_hd__clkbuf_1 _3073_ (.A(_1520_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _3074_ (.A0(net74),
    .A1(_1315_),
    .S(_1519_),
    .X(_1521_));
 sky130_fd_sc_hd__clkbuf_1 _3075_ (.A(_1521_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _3076_ (.A0(net151),
    .A1(_1317_),
    .S(_1519_),
    .X(_1522_));
 sky130_fd_sc_hd__clkbuf_1 _3077_ (.A(_1522_),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _3078_ (.A0(net350),
    .A1(_1319_),
    .S(_1519_),
    .X(_1523_));
 sky130_fd_sc_hd__clkbuf_1 _3079_ (.A(_1523_),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _3080_ (.A0(net246),
    .A1(_1321_),
    .S(_1519_),
    .X(_1524_));
 sky130_fd_sc_hd__clkbuf_1 _3081_ (.A(_1524_),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _3082_ (.A0(net156),
    .A1(_1323_),
    .S(_1519_),
    .X(_1525_));
 sky130_fd_sc_hd__clkbuf_1 _3083_ (.A(_1525_),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _3084_ (.A0(net279),
    .A1(_1325_),
    .S(_1519_),
    .X(_1526_));
 sky130_fd_sc_hd__clkbuf_1 _3085_ (.A(_1526_),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _3086_ (.A0(net267),
    .A1(_1327_),
    .S(_1519_),
    .X(_1527_));
 sky130_fd_sc_hd__clkbuf_1 _3087_ (.A(_1527_),
    .X(_0363_));
 sky130_fd_sc_hd__nand2_4 _3088_ (.A(_1451_),
    .B(_1509_),
    .Y(_1528_));
 sky130_fd_sc_hd__mux2_1 _3089_ (.A0(_1395_),
    .A1(\ram[50][0] ),
    .S(_1528_),
    .X(_1529_));
 sky130_fd_sc_hd__clkbuf_1 _3090_ (.A(_1529_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _3091_ (.A0(_1398_),
    .A1(\ram[50][1] ),
    .S(_1528_),
    .X(_1530_));
 sky130_fd_sc_hd__clkbuf_1 _3092_ (.A(_1530_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _3093_ (.A0(_1400_),
    .A1(\ram[50][2] ),
    .S(_1528_),
    .X(_1531_));
 sky130_fd_sc_hd__clkbuf_1 _3094_ (.A(_1531_),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_1 _3095_ (.A0(_1402_),
    .A1(\ram[50][3] ),
    .S(_1528_),
    .X(_1532_));
 sky130_fd_sc_hd__clkbuf_1 _3096_ (.A(_1532_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _3097_ (.A0(_1404_),
    .A1(\ram[50][4] ),
    .S(_1528_),
    .X(_1533_));
 sky130_fd_sc_hd__clkbuf_1 _3098_ (.A(_1533_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _3099_ (.A0(_1406_),
    .A1(\ram[50][5] ),
    .S(_1528_),
    .X(_1534_));
 sky130_fd_sc_hd__clkbuf_1 _3100_ (.A(_1534_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _3101_ (.A0(_1408_),
    .A1(net493),
    .S(_1528_),
    .X(_1535_));
 sky130_fd_sc_hd__clkbuf_1 _3102_ (.A(_1535_),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _3103_ (.A0(_1410_),
    .A1(net460),
    .S(_1528_),
    .X(_1536_));
 sky130_fd_sc_hd__clkbuf_1 _3104_ (.A(_1536_),
    .X(_0371_));
 sky130_fd_sc_hd__buf_2 _3105_ (.A(net7),
    .X(_1537_));
 sky130_fd_sc_hd__nand2_4 _3106_ (.A(_1127_),
    .B(_1509_),
    .Y(_1538_));
 sky130_fd_sc_hd__mux2_1 _3107_ (.A0(_1537_),
    .A1(net317),
    .S(_1538_),
    .X(_1539_));
 sky130_fd_sc_hd__clkbuf_1 _3108_ (.A(_1539_),
    .X(_0372_));
 sky130_fd_sc_hd__buf_2 _3109_ (.A(net8),
    .X(_1540_));
 sky130_fd_sc_hd__mux2_1 _3110_ (.A0(_1540_),
    .A1(net339),
    .S(_1538_),
    .X(_1541_));
 sky130_fd_sc_hd__clkbuf_1 _3111_ (.A(_1541_),
    .X(_0373_));
 sky130_fd_sc_hd__buf_2 _3112_ (.A(net9),
    .X(_1542_));
 sky130_fd_sc_hd__mux2_1 _3113_ (.A0(_1542_),
    .A1(net521),
    .S(_1538_),
    .X(_1543_));
 sky130_fd_sc_hd__clkbuf_1 _3114_ (.A(_1543_),
    .X(_0374_));
 sky130_fd_sc_hd__buf_2 _3115_ (.A(net10),
    .X(_1544_));
 sky130_fd_sc_hd__mux2_1 _3116_ (.A0(_1544_),
    .A1(net415),
    .S(_1538_),
    .X(_1545_));
 sky130_fd_sc_hd__clkbuf_1 _3117_ (.A(_1545_),
    .X(_0375_));
 sky130_fd_sc_hd__buf_2 _3118_ (.A(net11),
    .X(_1546_));
 sky130_fd_sc_hd__mux2_1 _3119_ (.A0(_1546_),
    .A1(net511),
    .S(_1538_),
    .X(_1547_));
 sky130_fd_sc_hd__clkbuf_1 _3120_ (.A(_1547_),
    .X(_0376_));
 sky130_fd_sc_hd__buf_2 _3121_ (.A(net12),
    .X(_1548_));
 sky130_fd_sc_hd__mux2_1 _3122_ (.A0(_1548_),
    .A1(net356),
    .S(_1538_),
    .X(_1549_));
 sky130_fd_sc_hd__clkbuf_1 _3123_ (.A(_1549_),
    .X(_0377_));
 sky130_fd_sc_hd__buf_2 _3124_ (.A(net13),
    .X(_1550_));
 sky130_fd_sc_hd__mux2_1 _3125_ (.A0(_1550_),
    .A1(net499),
    .S(_1538_),
    .X(_1551_));
 sky130_fd_sc_hd__clkbuf_1 _3126_ (.A(_1551_),
    .X(_0378_));
 sky130_fd_sc_hd__buf_2 _3127_ (.A(net14),
    .X(_1552_));
 sky130_fd_sc_hd__mux2_1 _3128_ (.A0(_1552_),
    .A1(net524),
    .S(_1538_),
    .X(_1553_));
 sky130_fd_sc_hd__clkbuf_1 _3129_ (.A(_1553_),
    .X(_0379_));
 sky130_fd_sc_hd__nand2_4 _3130_ (.A(_1470_),
    .B(_1509_),
    .Y(_1554_));
 sky130_fd_sc_hd__mux2_1 _3131_ (.A0(_1537_),
    .A1(net450),
    .S(_1554_),
    .X(_1555_));
 sky130_fd_sc_hd__clkbuf_1 _3132_ (.A(_1555_),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _3133_ (.A0(_1540_),
    .A1(net254),
    .S(_1554_),
    .X(_1556_));
 sky130_fd_sc_hd__clkbuf_1 _3134_ (.A(_1556_),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _3135_ (.A0(_1542_),
    .A1(net503),
    .S(_1554_),
    .X(_1557_));
 sky130_fd_sc_hd__clkbuf_1 _3136_ (.A(_1557_),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _3137_ (.A0(_1544_),
    .A1(net491),
    .S(_1554_),
    .X(_1558_));
 sky130_fd_sc_hd__clkbuf_1 _3138_ (.A(_1558_),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _3139_ (.A0(_1546_),
    .A1(net210),
    .S(_1554_),
    .X(_1559_));
 sky130_fd_sc_hd__clkbuf_1 _3140_ (.A(_1559_),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _3141_ (.A0(_1548_),
    .A1(net454),
    .S(_1554_),
    .X(_1560_));
 sky130_fd_sc_hd__clkbuf_1 _3142_ (.A(_1560_),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _3143_ (.A0(_1550_),
    .A1(net358),
    .S(_1554_),
    .X(_1561_));
 sky130_fd_sc_hd__clkbuf_1 _3144_ (.A(_1561_),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_1 _3145_ (.A0(_1552_),
    .A1(net429),
    .S(_1554_),
    .X(_1562_));
 sky130_fd_sc_hd__clkbuf_1 _3146_ (.A(_1562_),
    .X(_0387_));
 sky130_fd_sc_hd__nand2_4 _3147_ (.A(_1149_),
    .B(_1509_),
    .Y(_1563_));
 sky130_fd_sc_hd__mux2_1 _3148_ (.A0(_1537_),
    .A1(net225),
    .S(_1563_),
    .X(_1564_));
 sky130_fd_sc_hd__clkbuf_1 _3149_ (.A(_1564_),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _3150_ (.A0(_1540_),
    .A1(net361),
    .S(_1563_),
    .X(_1565_));
 sky130_fd_sc_hd__clkbuf_1 _3151_ (.A(_1565_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _3152_ (.A0(_1542_),
    .A1(net85),
    .S(_1563_),
    .X(_1566_));
 sky130_fd_sc_hd__clkbuf_1 _3153_ (.A(_1566_),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _3154_ (.A0(_1544_),
    .A1(net398),
    .S(_1563_),
    .X(_1567_));
 sky130_fd_sc_hd__clkbuf_1 _3155_ (.A(_1567_),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _3156_ (.A0(_1546_),
    .A1(net223),
    .S(_1563_),
    .X(_1568_));
 sky130_fd_sc_hd__clkbuf_1 _3157_ (.A(_1568_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _3158_ (.A0(_1548_),
    .A1(net414),
    .S(_1563_),
    .X(_1569_));
 sky130_fd_sc_hd__clkbuf_1 _3159_ (.A(_1569_),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _3160_ (.A0(_1550_),
    .A1(net461),
    .S(_1563_),
    .X(_1570_));
 sky130_fd_sc_hd__clkbuf_1 _3161_ (.A(_1570_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _3162_ (.A0(_1552_),
    .A1(net465),
    .S(_1563_),
    .X(_1571_));
 sky130_fd_sc_hd__clkbuf_1 _3163_ (.A(_1571_),
    .X(_0395_));
 sky130_fd_sc_hd__nand2_4 _3164_ (.A(_1161_),
    .B(_1509_),
    .Y(_1572_));
 sky130_fd_sc_hd__mux2_1 _3165_ (.A0(_1537_),
    .A1(net194),
    .S(_1572_),
    .X(_1573_));
 sky130_fd_sc_hd__clkbuf_1 _3166_ (.A(_1573_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _3167_ (.A0(_1540_),
    .A1(net269),
    .S(_1572_),
    .X(_1574_));
 sky130_fd_sc_hd__clkbuf_1 _3168_ (.A(_1574_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _3169_ (.A0(_1542_),
    .A1(net71),
    .S(_1572_),
    .X(_1575_));
 sky130_fd_sc_hd__clkbuf_1 _3170_ (.A(_1575_),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_1 _3171_ (.A0(_1544_),
    .A1(net432),
    .S(_1572_),
    .X(_1576_));
 sky130_fd_sc_hd__clkbuf_1 _3172_ (.A(_1576_),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _3173_ (.A0(_1546_),
    .A1(net229),
    .S(_1572_),
    .X(_1577_));
 sky130_fd_sc_hd__clkbuf_1 _3174_ (.A(_1577_),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _3175_ (.A0(_1548_),
    .A1(net431),
    .S(_1572_),
    .X(_1578_));
 sky130_fd_sc_hd__clkbuf_1 _3176_ (.A(_1578_),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _3177_ (.A0(_1550_),
    .A1(net315),
    .S(_1572_),
    .X(_1579_));
 sky130_fd_sc_hd__clkbuf_1 _3178_ (.A(_1579_),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _3179_ (.A0(_1552_),
    .A1(net294),
    .S(_1572_),
    .X(_1580_));
 sky130_fd_sc_hd__clkbuf_1 _3180_ (.A(_1580_),
    .X(_0403_));
 sky130_fd_sc_hd__nand2_4 _3181_ (.A(_1498_),
    .B(_1509_),
    .Y(_1581_));
 sky130_fd_sc_hd__mux2_1 _3182_ (.A0(_1537_),
    .A1(net405),
    .S(_1581_),
    .X(_1582_));
 sky130_fd_sc_hd__clkbuf_1 _3183_ (.A(_1582_),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_1 _3184_ (.A0(_1540_),
    .A1(net302),
    .S(_1581_),
    .X(_1583_));
 sky130_fd_sc_hd__clkbuf_1 _3185_ (.A(_1583_),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _3186_ (.A0(_1542_),
    .A1(net144),
    .S(_1581_),
    .X(_1584_));
 sky130_fd_sc_hd__clkbuf_1 _3187_ (.A(_1584_),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _3188_ (.A0(_1544_),
    .A1(net442),
    .S(_1581_),
    .X(_1585_));
 sky130_fd_sc_hd__clkbuf_1 _3189_ (.A(_1585_),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _3190_ (.A0(_1546_),
    .A1(net69),
    .S(_1581_),
    .X(_1586_));
 sky130_fd_sc_hd__clkbuf_1 _3191_ (.A(_1586_),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _3192_ (.A0(_1548_),
    .A1(net417),
    .S(_1581_),
    .X(_1587_));
 sky130_fd_sc_hd__clkbuf_1 _3193_ (.A(_1587_),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _3194_ (.A0(_1550_),
    .A1(net497),
    .S(_1581_),
    .X(_1588_));
 sky130_fd_sc_hd__clkbuf_1 _3195_ (.A(_1588_),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _3196_ (.A0(_1552_),
    .A1(net372),
    .S(_1581_),
    .X(_1589_));
 sky130_fd_sc_hd__clkbuf_1 _3197_ (.A(_1589_),
    .X(_0411_));
 sky130_fd_sc_hd__and3_1 _3198_ (.A(_0537_),
    .B(net5),
    .C(net6),
    .X(_1590_));
 sky130_fd_sc_hd__clkbuf_8 _3199_ (.A(_1590_),
    .X(_1591_));
 sky130_fd_sc_hd__nor2b_4 _3200_ (.A(_1094_),
    .B_N(_1591_),
    .Y(_1592_));
 sky130_fd_sc_hd__mux2_1 _3201_ (.A0(net325),
    .A1(_1312_),
    .S(_1592_),
    .X(_1593_));
 sky130_fd_sc_hd__clkbuf_1 _3202_ (.A(_1593_),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _3203_ (.A0(net408),
    .A1(_1315_),
    .S(_1592_),
    .X(_1594_));
 sky130_fd_sc_hd__clkbuf_1 _3204_ (.A(_1594_),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _3205_ (.A0(net30),
    .A1(_1317_),
    .S(_1592_),
    .X(_1595_));
 sky130_fd_sc_hd__clkbuf_1 _3206_ (.A(_1595_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _3207_ (.A0(net68),
    .A1(_1319_),
    .S(_1592_),
    .X(_1596_));
 sky130_fd_sc_hd__clkbuf_1 _3208_ (.A(_1596_),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _3209_ (.A0(net73),
    .A1(_1321_),
    .S(_1592_),
    .X(_1597_));
 sky130_fd_sc_hd__clkbuf_1 _3210_ (.A(_1597_),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _3211_ (.A0(net86),
    .A1(_1323_),
    .S(_1592_),
    .X(_1598_));
 sky130_fd_sc_hd__clkbuf_1 _3212_ (.A(_1598_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _3213_ (.A0(net367),
    .A1(_1325_),
    .S(_1592_),
    .X(_1599_));
 sky130_fd_sc_hd__clkbuf_1 _3214_ (.A(_1599_),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _3215_ (.A0(net108),
    .A1(_1327_),
    .S(_1592_),
    .X(_1600_));
 sky130_fd_sc_hd__clkbuf_1 _3216_ (.A(_1600_),
    .X(_0419_));
 sky130_fd_sc_hd__nand2_4 _3217_ (.A(_1441_),
    .B(_1591_),
    .Y(_1601_));
 sky130_fd_sc_hd__mux2_1 _3218_ (.A0(_1537_),
    .A1(net479),
    .S(_1601_),
    .X(_1602_));
 sky130_fd_sc_hd__clkbuf_1 _3219_ (.A(_1602_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _3220_ (.A0(_1540_),
    .A1(net467),
    .S(_1601_),
    .X(_1603_));
 sky130_fd_sc_hd__clkbuf_1 _3221_ (.A(_1603_),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _3222_ (.A0(_1542_),
    .A1(net240),
    .S(_1601_),
    .X(_1604_));
 sky130_fd_sc_hd__clkbuf_1 _3223_ (.A(_1604_),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _3224_ (.A0(_1544_),
    .A1(net80),
    .S(_1601_),
    .X(_1605_));
 sky130_fd_sc_hd__clkbuf_1 _3225_ (.A(_1605_),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _3226_ (.A0(_1546_),
    .A1(net228),
    .S(_1601_),
    .X(_1606_));
 sky130_fd_sc_hd__clkbuf_1 _3227_ (.A(_1606_),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _3228_ (.A0(_1548_),
    .A1(net173),
    .S(_1601_),
    .X(_1607_));
 sky130_fd_sc_hd__clkbuf_1 _3229_ (.A(_1607_),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _3230_ (.A0(_1550_),
    .A1(net35),
    .S(_1601_),
    .X(_1608_));
 sky130_fd_sc_hd__clkbuf_1 _3231_ (.A(_1608_),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _3232_ (.A0(_1552_),
    .A1(net334),
    .S(_1601_),
    .X(_1609_));
 sky130_fd_sc_hd__clkbuf_1 _3233_ (.A(_1609_),
    .X(_0427_));
 sky130_fd_sc_hd__nand2_4 _3234_ (.A(_1451_),
    .B(_1591_),
    .Y(_1610_));
 sky130_fd_sc_hd__mux2_1 _3235_ (.A0(_1537_),
    .A1(net423),
    .S(_1610_),
    .X(_1611_));
 sky130_fd_sc_hd__clkbuf_1 _3236_ (.A(_1611_),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _3237_ (.A0(_1540_),
    .A1(net480),
    .S(_1610_),
    .X(_1612_));
 sky130_fd_sc_hd__clkbuf_1 _3238_ (.A(_1612_),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _3239_ (.A0(_1542_),
    .A1(net250),
    .S(_1610_),
    .X(_1613_));
 sky130_fd_sc_hd__clkbuf_1 _3240_ (.A(_1613_),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _3241_ (.A0(_1544_),
    .A1(net168),
    .S(_1610_),
    .X(_1614_));
 sky130_fd_sc_hd__clkbuf_1 _3242_ (.A(_1614_),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _3243_ (.A0(_1546_),
    .A1(net131),
    .S(_1610_),
    .X(_1615_));
 sky130_fd_sc_hd__clkbuf_1 _3244_ (.A(_1615_),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _3245_ (.A0(_1548_),
    .A1(net79),
    .S(_1610_),
    .X(_1616_));
 sky130_fd_sc_hd__clkbuf_1 _3246_ (.A(_1616_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _3247_ (.A0(_1550_),
    .A1(net28),
    .S(_1610_),
    .X(_1617_));
 sky130_fd_sc_hd__clkbuf_1 _3248_ (.A(_1617_),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_1 _3249_ (.A0(_1552_),
    .A1(net278),
    .S(_1610_),
    .X(_1618_));
 sky130_fd_sc_hd__clkbuf_1 _3250_ (.A(_1618_),
    .X(_0435_));
 sky130_fd_sc_hd__nor2b_4 _3251_ (.A(_1053_),
    .B_N(_1072_),
    .Y(_1619_));
 sky130_fd_sc_hd__mux2_1 _3252_ (.A0(net133),
    .A1(net7),
    .S(_1619_),
    .X(_1620_));
 sky130_fd_sc_hd__clkbuf_1 _3253_ (.A(_1620_),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _3254_ (.A0(net154),
    .A1(net8),
    .S(_1619_),
    .X(_1621_));
 sky130_fd_sc_hd__clkbuf_1 _3255_ (.A(_1621_),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _3256_ (.A0(net227),
    .A1(net9),
    .S(_1619_),
    .X(_1622_));
 sky130_fd_sc_hd__clkbuf_1 _3257_ (.A(_1622_),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _3258_ (.A0(net298),
    .A1(net10),
    .S(_1619_),
    .X(_1623_));
 sky130_fd_sc_hd__clkbuf_1 _3259_ (.A(_1623_),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _3260_ (.A0(net283),
    .A1(net11),
    .S(_1619_),
    .X(_1624_));
 sky130_fd_sc_hd__clkbuf_1 _3261_ (.A(_1624_),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _3262_ (.A0(net182),
    .A1(net12),
    .S(_1619_),
    .X(_1625_));
 sky130_fd_sc_hd__clkbuf_1 _3263_ (.A(_1625_),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _3264_ (.A0(net436),
    .A1(net13),
    .S(_1619_),
    .X(_1626_));
 sky130_fd_sc_hd__clkbuf_1 _3265_ (.A(_1626_),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _3266_ (.A0(net420),
    .A1(net14),
    .S(_1619_),
    .X(_1627_));
 sky130_fd_sc_hd__clkbuf_1 _3267_ (.A(_1627_),
    .X(_0443_));
 sky130_fd_sc_hd__nand2_4 _3268_ (.A(_1470_),
    .B(_1591_),
    .Y(_1628_));
 sky130_fd_sc_hd__mux2_1 _3269_ (.A0(_1537_),
    .A1(net451),
    .S(_1628_),
    .X(_1629_));
 sky130_fd_sc_hd__clkbuf_1 _3270_ (.A(_1629_),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _3271_ (.A0(_1540_),
    .A1(net478),
    .S(_1628_),
    .X(_1630_));
 sky130_fd_sc_hd__clkbuf_1 _3272_ (.A(_1630_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _3273_ (.A0(_1542_),
    .A1(net103),
    .S(_1628_),
    .X(_1631_));
 sky130_fd_sc_hd__clkbuf_1 _3274_ (.A(_1631_),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_1 _3275_ (.A0(_1544_),
    .A1(net300),
    .S(_1628_),
    .X(_1632_));
 sky130_fd_sc_hd__clkbuf_1 _3276_ (.A(_1632_),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_1 _3277_ (.A0(_1546_),
    .A1(net492),
    .S(_1628_),
    .X(_1633_));
 sky130_fd_sc_hd__clkbuf_1 _3278_ (.A(_1633_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _3279_ (.A0(_1548_),
    .A1(net314),
    .S(_1628_),
    .X(_1634_));
 sky130_fd_sc_hd__clkbuf_1 _3280_ (.A(_1634_),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _3281_ (.A0(_1550_),
    .A1(net403),
    .S(_1628_),
    .X(_1635_));
 sky130_fd_sc_hd__clkbuf_1 _3282_ (.A(_1635_),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _3283_ (.A0(_1552_),
    .A1(net379),
    .S(_1628_),
    .X(_1636_));
 sky130_fd_sc_hd__clkbuf_1 _3284_ (.A(_1636_),
    .X(_0451_));
 sky130_fd_sc_hd__nand2_4 _3285_ (.A(_1149_),
    .B(_1591_),
    .Y(_1637_));
 sky130_fd_sc_hd__mux2_1 _3286_ (.A0(_1537_),
    .A1(net531),
    .S(_1637_),
    .X(_1638_));
 sky130_fd_sc_hd__clkbuf_1 _3287_ (.A(_1638_),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _3288_ (.A0(_1540_),
    .A1(\ram[61][1] ),
    .S(_1637_),
    .X(_1639_));
 sky130_fd_sc_hd__clkbuf_1 _3289_ (.A(_1639_),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _3290_ (.A0(_1542_),
    .A1(net424),
    .S(_1637_),
    .X(_1640_));
 sky130_fd_sc_hd__clkbuf_1 _3291_ (.A(_1640_),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _3292_ (.A0(_1544_),
    .A1(net459),
    .S(_1637_),
    .X(_1641_));
 sky130_fd_sc_hd__clkbuf_1 _3293_ (.A(_1641_),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _3294_ (.A0(_1546_),
    .A1(net439),
    .S(_1637_),
    .X(_1642_));
 sky130_fd_sc_hd__clkbuf_1 _3295_ (.A(_1642_),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_1 _3296_ (.A0(_1548_),
    .A1(net515),
    .S(_1637_),
    .X(_1643_));
 sky130_fd_sc_hd__clkbuf_1 _3297_ (.A(_1643_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _3298_ (.A0(_1550_),
    .A1(net255),
    .S(_1637_),
    .X(_1644_));
 sky130_fd_sc_hd__clkbuf_1 _3299_ (.A(_1644_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _3300_ (.A0(_1552_),
    .A1(net455),
    .S(_1637_),
    .X(_1645_));
 sky130_fd_sc_hd__clkbuf_1 _3301_ (.A(_1645_),
    .X(_0459_));
 sky130_fd_sc_hd__nand2_4 _3302_ (.A(_1161_),
    .B(_1591_),
    .Y(_1646_));
 sky130_fd_sc_hd__mux2_1 _3303_ (.A0(_1537_),
    .A1(net232),
    .S(_1646_),
    .X(_1647_));
 sky130_fd_sc_hd__clkbuf_1 _3304_ (.A(_1647_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _3305_ (.A0(_1540_),
    .A1(net53),
    .S(_1646_),
    .X(_1648_));
 sky130_fd_sc_hd__clkbuf_1 _3306_ (.A(_1648_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _3307_ (.A0(_1542_),
    .A1(net418),
    .S(_1646_),
    .X(_1649_));
 sky130_fd_sc_hd__clkbuf_1 _3308_ (.A(_1649_),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _3309_ (.A0(_1544_),
    .A1(net233),
    .S(_1646_),
    .X(_1650_));
 sky130_fd_sc_hd__clkbuf_1 _3310_ (.A(_1650_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _3311_ (.A0(_1546_),
    .A1(net235),
    .S(_1646_),
    .X(_1651_));
 sky130_fd_sc_hd__clkbuf_1 _3312_ (.A(_1651_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _3313_ (.A0(_1548_),
    .A1(net234),
    .S(_1646_),
    .X(_1652_));
 sky130_fd_sc_hd__clkbuf_1 _3314_ (.A(_1652_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _3315_ (.A0(_1550_),
    .A1(net411),
    .S(_1646_),
    .X(_1653_));
 sky130_fd_sc_hd__clkbuf_1 _3316_ (.A(_1653_),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _3317_ (.A0(_1552_),
    .A1(net438),
    .S(_1646_),
    .X(_1654_));
 sky130_fd_sc_hd__clkbuf_1 _3318_ (.A(_1654_),
    .X(_0467_));
 sky130_fd_sc_hd__nor2_4 _3319_ (.A(_1091_),
    .B(_1201_),
    .Y(_1655_));
 sky130_fd_sc_hd__mux2_1 _3320_ (.A0(net111),
    .A1(net7),
    .S(_1655_),
    .X(_1656_));
 sky130_fd_sc_hd__clkbuf_1 _3321_ (.A(_1656_),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _3322_ (.A0(net504),
    .A1(net8),
    .S(_1655_),
    .X(_1657_));
 sky130_fd_sc_hd__clkbuf_1 _3323_ (.A(_1657_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _3324_ (.A0(net231),
    .A1(net9),
    .S(_1655_),
    .X(_1658_));
 sky130_fd_sc_hd__clkbuf_1 _3325_ (.A(_1658_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _3326_ (.A0(net107),
    .A1(net10),
    .S(_1655_),
    .X(_1659_));
 sky130_fd_sc_hd__clkbuf_1 _3327_ (.A(_1659_),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _3328_ (.A0(net195),
    .A1(net11),
    .S(_1655_),
    .X(_1660_));
 sky130_fd_sc_hd__clkbuf_1 _3329_ (.A(_1660_),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _3330_ (.A0(net89),
    .A1(net12),
    .S(_1655_),
    .X(_1661_));
 sky130_fd_sc_hd__clkbuf_1 _3331_ (.A(_1661_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _3332_ (.A0(net243),
    .A1(net13),
    .S(_1655_),
    .X(_1662_));
 sky130_fd_sc_hd__clkbuf_1 _3333_ (.A(_1662_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _3334_ (.A0(net264),
    .A1(net14),
    .S(_1655_),
    .X(_1663_));
 sky130_fd_sc_hd__clkbuf_1 _3335_ (.A(_1663_),
    .X(_0475_));
 sky130_fd_sc_hd__nor2b_4 _3336_ (.A(_1053_),
    .B_N(_1159_),
    .Y(_1664_));
 sky130_fd_sc_hd__mux2_1 _3337_ (.A0(net175),
    .A1(net7),
    .S(_1664_),
    .X(_1665_));
 sky130_fd_sc_hd__clkbuf_1 _3338_ (.A(_1665_),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _3339_ (.A0(net44),
    .A1(net8),
    .S(_1664_),
    .X(_1666_));
 sky130_fd_sc_hd__clkbuf_1 _3340_ (.A(_1666_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _3341_ (.A0(net204),
    .A1(net9),
    .S(_1664_),
    .X(_1667_));
 sky130_fd_sc_hd__clkbuf_1 _3342_ (.A(_1667_),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _3343_ (.A0(net171),
    .A1(net10),
    .S(_1664_),
    .X(_1668_));
 sky130_fd_sc_hd__clkbuf_1 _3344_ (.A(_1668_),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _3345_ (.A0(net150),
    .A1(net11),
    .S(_1664_),
    .X(_1669_));
 sky130_fd_sc_hd__clkbuf_1 _3346_ (.A(_1669_),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _3347_ (.A0(net159),
    .A1(net12),
    .S(_1664_),
    .X(_1670_));
 sky130_fd_sc_hd__clkbuf_1 _3348_ (.A(_1670_),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _3349_ (.A0(net341),
    .A1(net13),
    .S(_1664_),
    .X(_1671_));
 sky130_fd_sc_hd__clkbuf_1 _3350_ (.A(_1671_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _3351_ (.A0(net208),
    .A1(net14),
    .S(_1664_),
    .X(_1672_));
 sky130_fd_sc_hd__clkbuf_1 _3352_ (.A(_1672_),
    .X(_0483_));
 sky130_fd_sc_hd__nand2_4 _3353_ (.A(_1498_),
    .B(_1591_),
    .Y(_1673_));
 sky130_fd_sc_hd__mux2_1 _3354_ (.A0(_1048_),
    .A1(net76),
    .S(_1673_),
    .X(_1674_));
 sky130_fd_sc_hd__clkbuf_1 _3355_ (.A(_1674_),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _3356_ (.A0(_1056_),
    .A1(net494),
    .S(_1673_),
    .X(_1675_));
 sky130_fd_sc_hd__clkbuf_1 _3357_ (.A(_1675_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _3358_ (.A0(_1058_),
    .A1(net124),
    .S(_1673_),
    .X(_1676_));
 sky130_fd_sc_hd__clkbuf_1 _3359_ (.A(_1676_),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _3360_ (.A0(_1060_),
    .A1(net458),
    .S(_1673_),
    .X(_1677_));
 sky130_fd_sc_hd__clkbuf_1 _3361_ (.A(_1677_),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _3362_ (.A0(_1062_),
    .A1(net364),
    .S(_1673_),
    .X(_1678_));
 sky130_fd_sc_hd__clkbuf_1 _3363_ (.A(_1678_),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _3364_ (.A0(_1064_),
    .A1(net147),
    .S(_1673_),
    .X(_1679_));
 sky130_fd_sc_hd__clkbuf_1 _3365_ (.A(_1679_),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _3366_ (.A0(_1066_),
    .A1(net366),
    .S(_1673_),
    .X(_1680_));
 sky130_fd_sc_hd__clkbuf_1 _3367_ (.A(_1680_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _3368_ (.A0(_1068_),
    .A1(net396),
    .S(_1673_),
    .X(_1681_));
 sky130_fd_sc_hd__clkbuf_1 _3369_ (.A(_1681_),
    .X(_0491_));
 sky130_fd_sc_hd__nand2_4 _3370_ (.A(_1127_),
    .B(_1591_),
    .Y(_1682_));
 sky130_fd_sc_hd__mux2_1 _3371_ (.A0(_1048_),
    .A1(net188),
    .S(_1682_),
    .X(_1683_));
 sky130_fd_sc_hd__clkbuf_1 _3372_ (.A(_1683_),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _3373_ (.A0(_1056_),
    .A1(net397),
    .S(_1682_),
    .X(_1684_));
 sky130_fd_sc_hd__clkbuf_1 _3374_ (.A(_1684_),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _3375_ (.A0(_1058_),
    .A1(net290),
    .S(_1682_),
    .X(_1685_));
 sky130_fd_sc_hd__clkbuf_1 _3376_ (.A(_1685_),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _3377_ (.A0(_1060_),
    .A1(net306),
    .S(_1682_),
    .X(_1686_));
 sky130_fd_sc_hd__clkbuf_1 _3378_ (.A(_1686_),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_1 _3379_ (.A0(_1062_),
    .A1(net193),
    .S(_1682_),
    .X(_1687_));
 sky130_fd_sc_hd__clkbuf_1 _3380_ (.A(_1687_),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _3381_ (.A0(_1064_),
    .A1(net413),
    .S(_1682_),
    .X(_1688_));
 sky130_fd_sc_hd__clkbuf_1 _3382_ (.A(_1688_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _3383_ (.A0(_1066_),
    .A1(net57),
    .S(_1682_),
    .X(_1689_));
 sky130_fd_sc_hd__clkbuf_1 _3384_ (.A(_1689_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _3385_ (.A0(_1068_),
    .A1(net342),
    .S(_1682_),
    .X(_1690_));
 sky130_fd_sc_hd__clkbuf_1 _3386_ (.A(_1690_),
    .X(_0499_));
 sky130_fd_sc_hd__nand2_4 _3387_ (.A(_1441_),
    .B(_1509_),
    .Y(_1691_));
 sky130_fd_sc_hd__mux2_1 _3388_ (.A0(_1048_),
    .A1(net447),
    .S(_1691_),
    .X(_1692_));
 sky130_fd_sc_hd__clkbuf_1 _3389_ (.A(_1692_),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _3390_ (.A0(_1056_),
    .A1(net400),
    .S(_1691_),
    .X(_1693_));
 sky130_fd_sc_hd__clkbuf_1 _3391_ (.A(_1693_),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _3392_ (.A0(_1058_),
    .A1(net529),
    .S(_1691_),
    .X(_1694_));
 sky130_fd_sc_hd__clkbuf_1 _3393_ (.A(_1694_),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _3394_ (.A0(_1060_),
    .A1(net496),
    .S(_1691_),
    .X(_1695_));
 sky130_fd_sc_hd__clkbuf_1 _3395_ (.A(_1695_),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_1 _3396_ (.A0(_1062_),
    .A1(net416),
    .S(_1691_),
    .X(_1696_));
 sky130_fd_sc_hd__clkbuf_1 _3397_ (.A(_1696_),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_1 _3398_ (.A0(_1064_),
    .A1(net362),
    .S(_1691_),
    .X(_1697_));
 sky130_fd_sc_hd__clkbuf_1 _3399_ (.A(_1697_),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _3400_ (.A0(_1066_),
    .A1(net483),
    .S(_1691_),
    .X(_1698_));
 sky130_fd_sc_hd__clkbuf_1 _3401_ (.A(_1698_),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _3402_ (.A0(_1068_),
    .A1(net46),
    .S(_1691_),
    .X(_1699_));
 sky130_fd_sc_hd__clkbuf_1 _3403_ (.A(_1699_),
    .X(_0507_));
 sky130_fd_sc_hd__nand2_4 _3404_ (.A(_1127_),
    .B(_1238_),
    .Y(_1700_));
 sky130_fd_sc_hd__mux2_1 _3405_ (.A0(_1048_),
    .A1(net441),
    .S(_1700_),
    .X(_1701_));
 sky130_fd_sc_hd__clkbuf_1 _3406_ (.A(_1701_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _3407_ (.A0(_1056_),
    .A1(net374),
    .S(_1700_),
    .X(_1702_));
 sky130_fd_sc_hd__clkbuf_1 _3408_ (.A(_1702_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _3409_ (.A0(_1058_),
    .A1(net296),
    .S(_1700_),
    .X(_1703_));
 sky130_fd_sc_hd__clkbuf_1 _3410_ (.A(_1703_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _3411_ (.A0(_1060_),
    .A1(net181),
    .S(_1700_),
    .X(_1704_));
 sky130_fd_sc_hd__clkbuf_1 _3412_ (.A(_1704_),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _3413_ (.A0(_1062_),
    .A1(net281),
    .S(_1700_),
    .X(_1705_));
 sky130_fd_sc_hd__clkbuf_1 _3414_ (.A(_1705_),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _3415_ (.A0(_1064_),
    .A1(net527),
    .S(_1700_),
    .X(_1706_));
 sky130_fd_sc_hd__clkbuf_1 _3416_ (.A(_1706_),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _3417_ (.A0(_1066_),
    .A1(net399),
    .S(_1700_),
    .X(_1707_));
 sky130_fd_sc_hd__clkbuf_1 _3418_ (.A(_1707_),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _3419_ (.A0(_1068_),
    .A1(net98),
    .S(_1700_),
    .X(_1708_));
 sky130_fd_sc_hd__clkbuf_1 _3420_ (.A(_1708_),
    .X(_0515_));
 sky130_fd_sc_hd__nor2_4 _3421_ (.A(_1171_),
    .B(_1348_),
    .Y(_1709_));
 sky130_fd_sc_hd__mux2_1 _3422_ (.A0(net401),
    .A1(net7),
    .S(_1709_),
    .X(_1710_));
 sky130_fd_sc_hd__clkbuf_1 _3423_ (.A(_1710_),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _3424_ (.A0(net388),
    .A1(net8),
    .S(_1709_),
    .X(_1711_));
 sky130_fd_sc_hd__clkbuf_1 _3425_ (.A(_1711_),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _3426_ (.A0(net344),
    .A1(net9),
    .S(_1709_),
    .X(_1712_));
 sky130_fd_sc_hd__clkbuf_1 _3427_ (.A(_1712_),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_1 _3428_ (.A0(net286),
    .A1(net10),
    .S(_1709_),
    .X(_1713_));
 sky130_fd_sc_hd__clkbuf_1 _3429_ (.A(_1713_),
    .X(_0519_));
 sky130_fd_sc_hd__mux2_1 _3430_ (.A0(net191),
    .A1(net11),
    .S(_1709_),
    .X(_1714_));
 sky130_fd_sc_hd__clkbuf_1 _3431_ (.A(_1714_),
    .X(_0520_));
 sky130_fd_sc_hd__mux2_1 _3432_ (.A0(net310),
    .A1(net12),
    .S(_1709_),
    .X(_1715_));
 sky130_fd_sc_hd__clkbuf_1 _3433_ (.A(_1715_),
    .X(_0521_));
 sky130_fd_sc_hd__mux2_1 _3434_ (.A0(net33),
    .A1(net13),
    .S(_1709_),
    .X(_1716_));
 sky130_fd_sc_hd__clkbuf_1 _3435_ (.A(_1716_),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_1 _3436_ (.A0(net332),
    .A1(net14),
    .S(_1709_),
    .X(_1717_));
 sky130_fd_sc_hd__clkbuf_1 _3437_ (.A(_1717_),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_1 _3438_ (.A0(_0530_),
    .A1(net463),
    .S(_0531_),
    .X(_1718_));
 sky130_fd_sc_hd__clkbuf_1 _3439_ (.A(_1718_),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_1 _3440_ (.A0(_0533_),
    .A1(net385),
    .S(_0531_),
    .X(_1719_));
 sky130_fd_sc_hd__clkbuf_1 _3441_ (.A(_1719_),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_1 _3442_ (.A0(_0535_),
    .A1(net476),
    .S(_0531_),
    .X(_1720_));
 sky130_fd_sc_hd__clkbuf_1 _3443_ (.A(_1720_),
    .X(_0526_));
 sky130_fd_sc_hd__mux2_1 _3444_ (.A0(_0537_),
    .A1(net197),
    .S(_0531_),
    .X(_1721_));
 sky130_fd_sc_hd__clkbuf_1 _3445_ (.A(_1721_),
    .X(_0527_));
 sky130_fd_sc_hd__mux2_1 _3446_ (.A0(net5),
    .A1(net282),
    .S(net15),
    .X(_1722_));
 sky130_fd_sc_hd__clkbuf_1 _3447_ (.A(_1722_),
    .X(_0528_));
 sky130_fd_sc_hd__mux2_1 _3448_ (.A0(_0540_),
    .A1(net24),
    .S(net15),
    .X(_1723_));
 sky130_fd_sc_hd__clkbuf_1 _3449_ (.A(_1723_),
    .X(_0529_));
 sky130_fd_sc_hd__dfxtp_1 _3450_ (.CLK(clknet_leaf_39_clk),
    .D(_0012_),
    .Q(\ram[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3451_ (.CLK(clknet_leaf_39_clk),
    .D(_0013_),
    .Q(\ram[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3452_ (.CLK(clknet_leaf_41_clk),
    .D(_0014_),
    .Q(\ram[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3453_ (.CLK(clknet_leaf_40_clk),
    .D(_0015_),
    .Q(\ram[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3454_ (.CLK(clknet_leaf_40_clk),
    .D(_0016_),
    .Q(\ram[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3455_ (.CLK(clknet_leaf_39_clk),
    .D(_0017_),
    .Q(\ram[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3456_ (.CLK(clknet_leaf_37_clk),
    .D(_0018_),
    .Q(\ram[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3457_ (.CLK(clknet_leaf_37_clk),
    .D(_0019_),
    .Q(\ram[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3458_ (.CLK(clknet_leaf_8_clk),
    .D(_0020_),
    .Q(\ram[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3459_ (.CLK(clknet_leaf_0_clk),
    .D(_0021_),
    .Q(\ram[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3460_ (.CLK(clknet_leaf_6_clk),
    .D(_0022_),
    .Q(\ram[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3461_ (.CLK(clknet_leaf_7_clk),
    .D(_0023_),
    .Q(\ram[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3462_ (.CLK(clknet_leaf_7_clk),
    .D(_0024_),
    .Q(\ram[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3463_ (.CLK(clknet_leaf_1_clk),
    .D(_0025_),
    .Q(\ram[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3464_ (.CLK(clknet_leaf_2_clk),
    .D(_0026_),
    .Q(\ram[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3465_ (.CLK(clknet_leaf_3_clk),
    .D(_0027_),
    .Q(\ram[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3466_ (.CLK(clknet_leaf_5_clk),
    .D(_0028_),
    .Q(\ram[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3467_ (.CLK(clknet_leaf_10_clk),
    .D(_0029_),
    .Q(\ram[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3468_ (.CLK(clknet_leaf_10_clk),
    .D(_0030_),
    .Q(\ram[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3469_ (.CLK(clknet_leaf_12_clk),
    .D(_0031_),
    .Q(\ram[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3470_ (.CLK(clknet_leaf_10_clk),
    .D(_0032_),
    .Q(\ram[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3471_ (.CLK(clknet_leaf_5_clk),
    .D(_0033_),
    .Q(\ram[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3472_ (.CLK(clknet_leaf_13_clk),
    .D(_0034_),
    .Q(\ram[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3473_ (.CLK(clknet_leaf_13_clk),
    .D(_0035_),
    .Q(\ram[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3474_ (.CLK(clknet_leaf_42_clk),
    .D(_0036_),
    .Q(\ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3475_ (.CLK(clknet_leaf_39_clk),
    .D(_0037_),
    .Q(\ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3476_ (.CLK(clknet_leaf_41_clk),
    .D(_0038_),
    .Q(\ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3477_ (.CLK(clknet_leaf_34_clk),
    .D(_0039_),
    .Q(\ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3478_ (.CLK(clknet_leaf_41_clk),
    .D(_0040_),
    .Q(\ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3479_ (.CLK(clknet_leaf_40_clk),
    .D(_0041_),
    .Q(\ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3480_ (.CLK(clknet_leaf_36_clk),
    .D(_0042_),
    .Q(\ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3481_ (.CLK(clknet_leaf_36_clk),
    .D(_0043_),
    .Q(\ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3482_ (.CLK(clknet_leaf_10_clk),
    .D(_0044_),
    .Q(\ram[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3483_ (.CLK(clknet_leaf_10_clk),
    .D(_0045_),
    .Q(\ram[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3484_ (.CLK(clknet_leaf_10_clk),
    .D(_0046_),
    .Q(\ram[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3485_ (.CLK(clknet_leaf_11_clk),
    .D(_0047_),
    .Q(\ram[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3486_ (.CLK(clknet_leaf_10_clk),
    .D(_0048_),
    .Q(\ram[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3487_ (.CLK(clknet_leaf_5_clk),
    .D(_0049_),
    .Q(\ram[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3488_ (.CLK(clknet_leaf_13_clk),
    .D(_0050_),
    .Q(\ram[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3489_ (.CLK(clknet_leaf_13_clk),
    .D(_0051_),
    .Q(\ram[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3490_ (.CLK(clknet_leaf_10_clk),
    .D(_0052_),
    .Q(\ram[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3491_ (.CLK(clknet_leaf_10_clk),
    .D(_0053_),
    .Q(\ram[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3492_ (.CLK(clknet_leaf_10_clk),
    .D(_0054_),
    .Q(\ram[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3493_ (.CLK(clknet_leaf_11_clk),
    .D(_0055_),
    .Q(\ram[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3494_ (.CLK(clknet_leaf_10_clk),
    .D(_0056_),
    .Q(\ram[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3495_ (.CLK(clknet_leaf_5_clk),
    .D(_0057_),
    .Q(\ram[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3496_ (.CLK(clknet_leaf_13_clk),
    .D(_0058_),
    .Q(\ram[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3497_ (.CLK(clknet_leaf_12_clk),
    .D(_0059_),
    .Q(\ram[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3498_ (.CLK(clknet_leaf_8_clk),
    .D(_0060_),
    .Q(\ram[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3499_ (.CLK(clknet_leaf_9_clk),
    .D(_0061_),
    .Q(\ram[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3500_ (.CLK(clknet_leaf_9_clk),
    .D(_0062_),
    .Q(\ram[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3501_ (.CLK(clknet_leaf_10_clk),
    .D(_0063_),
    .Q(\ram[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3502_ (.CLK(clknet_leaf_10_clk),
    .D(_0064_),
    .Q(\ram[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3503_ (.CLK(clknet_leaf_8_clk),
    .D(_0065_),
    .Q(\ram[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3504_ (.CLK(clknet_leaf_13_clk),
    .D(_0066_),
    .Q(\ram[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3505_ (.CLK(clknet_leaf_13_clk),
    .D(_0067_),
    .Q(\ram[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3506_ (.CLK(clknet_leaf_8_clk),
    .D(_0068_),
    .Q(\ram[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3507_ (.CLK(clknet_leaf_9_clk),
    .D(_0069_),
    .Q(\ram[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3508_ (.CLK(clknet_leaf_9_clk),
    .D(_0070_),
    .Q(\ram[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3509_ (.CLK(clknet_leaf_10_clk),
    .D(_0071_),
    .Q(\ram[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3510_ (.CLK(clknet_leaf_8_clk),
    .D(_0072_),
    .Q(\ram[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3511_ (.CLK(clknet_leaf_8_clk),
    .D(_0073_),
    .Q(\ram[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3512_ (.CLK(clknet_leaf_13_clk),
    .D(_0074_),
    .Q(\ram[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3513_ (.CLK(clknet_leaf_13_clk),
    .D(_0075_),
    .Q(\ram[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3514_ (.CLK(clknet_leaf_8_clk),
    .D(_0076_),
    .Q(\ram[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3515_ (.CLK(clknet_leaf_9_clk),
    .D(_0077_),
    .Q(\ram[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3516_ (.CLK(clknet_leaf_9_clk),
    .D(_0078_),
    .Q(\ram[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3517_ (.CLK(clknet_leaf_10_clk),
    .D(_0079_),
    .Q(\ram[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3518_ (.CLK(clknet_leaf_9_clk),
    .D(_0080_),
    .Q(\ram[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3519_ (.CLK(clknet_leaf_8_clk),
    .D(_0081_),
    .Q(\ram[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3520_ (.CLK(clknet_leaf_4_clk),
    .D(_0082_),
    .Q(\ram[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3521_ (.CLK(clknet_leaf_13_clk),
    .D(_0083_),
    .Q(\ram[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3522_ (.CLK(clknet_leaf_8_clk),
    .D(_0084_),
    .Q(\ram[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3523_ (.CLK(clknet_leaf_9_clk),
    .D(_0085_),
    .Q(\ram[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3524_ (.CLK(clknet_leaf_9_clk),
    .D(_0086_),
    .Q(\ram[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3525_ (.CLK(clknet_leaf_10_clk),
    .D(_0087_),
    .Q(\ram[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3526_ (.CLK(clknet_leaf_8_clk),
    .D(_0088_),
    .Q(\ram[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3527_ (.CLK(clknet_leaf_8_clk),
    .D(_0089_),
    .Q(\ram[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3528_ (.CLK(clknet_leaf_4_clk),
    .D(_0090_),
    .Q(\ram[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3529_ (.CLK(clknet_leaf_13_clk),
    .D(_0091_),
    .Q(\ram[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3530_ (.CLK(clknet_leaf_43_clk),
    .D(_0092_),
    .Q(\ram[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3531_ (.CLK(clknet_leaf_44_clk),
    .D(_0093_),
    .Q(\ram[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3532_ (.CLK(clknet_leaf_42_clk),
    .D(_0094_),
    .Q(\ram[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3533_ (.CLK(clknet_leaf_42_clk),
    .D(_0095_),
    .Q(\ram[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3534_ (.CLK(clknet_leaf_43_clk),
    .D(_0096_),
    .Q(\ram[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3535_ (.CLK(clknet_leaf_44_clk),
    .D(_0097_),
    .Q(\ram[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3536_ (.CLK(clknet_leaf_38_clk),
    .D(_0098_),
    .Q(\ram[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3537_ (.CLK(clknet_leaf_38_clk),
    .D(_0099_),
    .Q(\ram[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3538_ (.CLK(clknet_leaf_43_clk),
    .D(_0100_),
    .Q(\ram[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3539_ (.CLK(clknet_leaf_44_clk),
    .D(_0101_),
    .Q(\ram[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3540_ (.CLK(clknet_leaf_42_clk),
    .D(_0102_),
    .Q(\ram[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3541_ (.CLK(clknet_leaf_41_clk),
    .D(_0103_),
    .Q(\ram[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3542_ (.CLK(clknet_leaf_43_clk),
    .D(_0104_),
    .Q(\ram[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3543_ (.CLK(clknet_leaf_2_clk),
    .D(_0105_),
    .Q(\ram[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3544_ (.CLK(clknet_leaf_38_clk),
    .D(_0106_),
    .Q(\ram[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3545_ (.CLK(clknet_leaf_38_clk),
    .D(_0107_),
    .Q(\ram[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3546_ (.CLK(clknet_leaf_43_clk),
    .D(_0108_),
    .Q(\ram[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3547_ (.CLK(clknet_leaf_44_clk),
    .D(_0109_),
    .Q(\ram[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3548_ (.CLK(clknet_leaf_43_clk),
    .D(_0110_),
    .Q(\ram[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3549_ (.CLK(clknet_leaf_43_clk),
    .D(_0111_),
    .Q(\ram[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3550_ (.CLK(clknet_leaf_43_clk),
    .D(_0112_),
    .Q(\ram[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3551_ (.CLK(clknet_leaf_44_clk),
    .D(_0113_),
    .Q(\ram[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3552_ (.CLK(clknet_leaf_39_clk),
    .D(_0114_),
    .Q(\ram[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3553_ (.CLK(clknet_leaf_38_clk),
    .D(_0115_),
    .Q(\ram[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3554_ (.CLK(clknet_leaf_42_clk),
    .D(_0116_),
    .Q(\ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3555_ (.CLK(clknet_leaf_2_clk),
    .D(_0117_),
    .Q(\ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3556_ (.CLK(clknet_leaf_41_clk),
    .D(_0118_),
    .Q(\ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3557_ (.CLK(clknet_leaf_40_clk),
    .D(_0119_),
    .Q(\ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3558_ (.CLK(clknet_leaf_41_clk),
    .D(_0120_),
    .Q(\ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3559_ (.CLK(clknet_leaf_40_clk),
    .D(_0121_),
    .Q(\ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3560_ (.CLK(clknet_leaf_39_clk),
    .D(_0122_),
    .Q(\ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3561_ (.CLK(clknet_leaf_37_clk),
    .D(_0123_),
    .Q(\ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3562_ (.CLK(clknet_leaf_6_clk),
    .D(_0124_),
    .Q(\ram[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3563_ (.CLK(clknet_leaf_1_clk),
    .D(_0125_),
    .Q(\ram[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3564_ (.CLK(clknet_leaf_6_clk),
    .D(_0126_),
    .Q(\ram[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3565_ (.CLK(clknet_leaf_6_clk),
    .D(_0127_),
    .Q(\ram[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3566_ (.CLK(clknet_leaf_6_clk),
    .D(_0128_),
    .Q(\ram[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3567_ (.CLK(clknet_leaf_1_clk),
    .D(_0129_),
    .Q(\ram[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3568_ (.CLK(clknet_leaf_3_clk),
    .D(_0130_),
    .Q(\ram[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3569_ (.CLK(clknet_leaf_3_clk),
    .D(_0131_),
    .Q(\ram[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3570_ (.CLK(clknet_leaf_6_clk),
    .D(_0132_),
    .Q(\ram[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3571_ (.CLK(clknet_leaf_1_clk),
    .D(_0133_),
    .Q(\ram[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3572_ (.CLK(clknet_leaf_6_clk),
    .D(_0134_),
    .Q(\ram[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3573_ (.CLK(clknet_leaf_6_clk),
    .D(_0135_),
    .Q(\ram[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3574_ (.CLK(clknet_leaf_6_clk),
    .D(_0136_),
    .Q(\ram[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3575_ (.CLK(clknet_leaf_1_clk),
    .D(_0137_),
    .Q(\ram[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3576_ (.CLK(clknet_leaf_3_clk),
    .D(_0138_),
    .Q(\ram[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3577_ (.CLK(clknet_leaf_3_clk),
    .D(_0139_),
    .Q(\ram[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3578_ (.CLK(clknet_leaf_4_clk),
    .D(_0140_),
    .Q(\ram[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3579_ (.CLK(clknet_leaf_2_clk),
    .D(_0141_),
    .Q(\ram[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3580_ (.CLK(clknet_leaf_5_clk),
    .D(_0142_),
    .Q(\ram[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3581_ (.CLK(clknet_leaf_5_clk),
    .D(_0143_),
    .Q(\ram[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3582_ (.CLK(clknet_leaf_5_clk),
    .D(_0144_),
    .Q(\ram[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3583_ (.CLK(clknet_leaf_1_clk),
    .D(_0145_),
    .Q(\ram[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3584_ (.CLK(clknet_leaf_3_clk),
    .D(_0146_),
    .Q(\ram[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3585_ (.CLK(clknet_leaf_4_clk),
    .D(_0147_),
    .Q(\ram[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3586_ (.CLK(clknet_leaf_4_clk),
    .D(_0148_),
    .Q(\ram[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3587_ (.CLK(clknet_leaf_2_clk),
    .D(_0149_),
    .Q(\ram[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3588_ (.CLK(clknet_leaf_4_clk),
    .D(_0150_),
    .Q(\ram[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3589_ (.CLK(clknet_leaf_5_clk),
    .D(_0151_),
    .Q(\ram[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3590_ (.CLK(clknet_leaf_5_clk),
    .D(_0152_),
    .Q(\ram[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3591_ (.CLK(clknet_leaf_1_clk),
    .D(_0153_),
    .Q(\ram[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3592_ (.CLK(clknet_leaf_2_clk),
    .D(_0154_),
    .Q(\ram[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3593_ (.CLK(clknet_leaf_4_clk),
    .D(_0155_),
    .Q(\ram[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3594_ (.CLK(clknet_leaf_2_clk),
    .D(_0156_),
    .Q(\ram[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3595_ (.CLK(clknet_leaf_44_clk),
    .D(_0157_),
    .Q(\ram[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3596_ (.CLK(clknet_leaf_44_clk),
    .D(_0158_),
    .Q(\ram[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3597_ (.CLK(clknet_leaf_44_clk),
    .D(_0159_),
    .Q(\ram[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3598_ (.CLK(clknet_leaf_0_clk),
    .D(_0160_),
    .Q(\ram[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3599_ (.CLK(clknet_leaf_1_clk),
    .D(_0161_),
    .Q(\ram[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3600_ (.CLK(clknet_leaf_38_clk),
    .D(_0162_),
    .Q(\ram[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3601_ (.CLK(clknet_leaf_37_clk),
    .D(_0163_),
    .Q(\ram[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3602_ (.CLK(clknet_leaf_2_clk),
    .D(_0164_),
    .Q(\ram[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3603_ (.CLK(clknet_leaf_1_clk),
    .D(_0165_),
    .Q(\ram[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3604_ (.CLK(clknet_leaf_44_clk),
    .D(_0166_),
    .Q(\ram[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3605_ (.CLK(clknet_leaf_44_clk),
    .D(_0167_),
    .Q(\ram[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3606_ (.CLK(clknet_leaf_1_clk),
    .D(_0168_),
    .Q(\ram[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3607_ (.CLK(clknet_leaf_44_clk),
    .D(_0169_),
    .Q(\ram[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3608_ (.CLK(clknet_leaf_2_clk),
    .D(_0170_),
    .Q(\ram[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3609_ (.CLK(clknet_leaf_38_clk),
    .D(_0171_),
    .Q(\ram[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3610_ (.CLK(clknet_leaf_1_clk),
    .D(_0172_),
    .Q(\ram[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3611_ (.CLK(clknet_leaf_0_clk),
    .D(_0173_),
    .Q(\ram[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3612_ (.CLK(clknet_leaf_0_clk),
    .D(_0174_),
    .Q(\ram[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3613_ (.CLK(clknet_leaf_0_clk),
    .D(_0175_),
    .Q(\ram[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3614_ (.CLK(clknet_leaf_0_clk),
    .D(_0176_),
    .Q(\ram[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3615_ (.CLK(clknet_leaf_44_clk),
    .D(_0177_),
    .Q(\ram[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3616_ (.CLK(clknet_leaf_2_clk),
    .D(_0178_),
    .Q(\ram[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3617_ (.CLK(clknet_leaf_2_clk),
    .D(_0179_),
    .Q(\ram[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3618_ (.CLK(clknet_leaf_1_clk),
    .D(_0180_),
    .Q(\ram[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3619_ (.CLK(clknet_leaf_0_clk),
    .D(_0181_),
    .Q(\ram[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3620_ (.CLK(clknet_leaf_0_clk),
    .D(_0182_),
    .Q(\ram[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3621_ (.CLK(clknet_leaf_0_clk),
    .D(_0183_),
    .Q(\ram[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3622_ (.CLK(clknet_leaf_0_clk),
    .D(_0184_),
    .Q(\ram[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3623_ (.CLK(clknet_leaf_1_clk),
    .D(_0185_),
    .Q(\ram[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3624_ (.CLK(clknet_leaf_2_clk),
    .D(_0186_),
    .Q(\ram[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3625_ (.CLK(clknet_leaf_2_clk),
    .D(_0187_),
    .Q(\ram[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3626_ (.CLK(clknet_leaf_5_clk),
    .D(_0188_),
    .Q(\ram[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3627_ (.CLK(clknet_leaf_0_clk),
    .D(_0189_),
    .Q(\ram[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3628_ (.CLK(clknet_leaf_6_clk),
    .D(_0190_),
    .Q(\ram[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3629_ (.CLK(clknet_leaf_7_clk),
    .D(_0191_),
    .Q(\ram[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3630_ (.CLK(clknet_leaf_7_clk),
    .D(_0192_),
    .Q(\ram[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3631_ (.CLK(clknet_leaf_1_clk),
    .D(_0193_),
    .Q(\ram[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3632_ (.CLK(clknet_leaf_2_clk),
    .D(_0194_),
    .Q(\ram[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3633_ (.CLK(clknet_leaf_3_clk),
    .D(_0195_),
    .Q(\ram[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3634_ (.CLK(clknet_leaf_42_clk),
    .D(_0196_),
    .Q(\ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3635_ (.CLK(clknet_leaf_42_clk),
    .D(_0197_),
    .Q(\ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3636_ (.CLK(clknet_leaf_42_clk),
    .D(_0198_),
    .Q(\ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3637_ (.CLK(clknet_leaf_40_clk),
    .D(_0199_),
    .Q(\ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3638_ (.CLK(clknet_leaf_41_clk),
    .D(_0200_),
    .Q(\ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3639_ (.CLK(clknet_leaf_41_clk),
    .D(_0201_),
    .Q(\ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3640_ (.CLK(clknet_leaf_35_clk),
    .D(_0202_),
    .Q(\ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3641_ (.CLK(clknet_leaf_37_clk),
    .D(_0203_),
    .Q(\ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3642_ (.CLK(clknet_leaf_7_clk),
    .D(_0204_),
    .Q(\ram[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3643_ (.CLK(clknet_leaf_0_clk),
    .D(_0205_),
    .Q(\ram[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3644_ (.CLK(clknet_leaf_7_clk),
    .D(_0206_),
    .Q(\ram[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3645_ (.CLK(clknet_leaf_7_clk),
    .D(_0207_),
    .Q(\ram[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3646_ (.CLK(clknet_leaf_7_clk),
    .D(_0208_),
    .Q(\ram[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3647_ (.CLK(clknet_leaf_8_clk),
    .D(_0209_),
    .Q(\ram[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3648_ (.CLK(clknet_leaf_3_clk),
    .D(_0210_),
    .Q(\ram[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3649_ (.CLK(clknet_leaf_14_clk),
    .D(_0211_),
    .Q(\ram[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3650_ (.CLK(clknet_leaf_8_clk),
    .D(_0212_),
    .Q(\ram[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3651_ (.CLK(clknet_leaf_0_clk),
    .D(_0213_),
    .Q(\ram[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3652_ (.CLK(clknet_leaf_7_clk),
    .D(_0214_),
    .Q(\ram[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3653_ (.CLK(clknet_leaf_7_clk),
    .D(_0215_),
    .Q(\ram[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3654_ (.CLK(clknet_leaf_7_clk),
    .D(_0216_),
    .Q(\ram[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3655_ (.CLK(clknet_leaf_8_clk),
    .D(_0217_),
    .Q(\ram[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3656_ (.CLK(clknet_leaf_3_clk),
    .D(_0218_),
    .Q(\ram[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3657_ (.CLK(clknet_leaf_3_clk),
    .D(_0219_),
    .Q(\ram[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3658_ (.CLK(clknet_leaf_16_clk),
    .D(_0220_),
    .Q(\ram[32][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3659_ (.CLK(clknet_leaf_17_clk),
    .D(_0221_),
    .Q(\ram[32][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3660_ (.CLK(clknet_leaf_11_clk),
    .D(_0222_),
    .Q(\ram[32][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3661_ (.CLK(clknet_leaf_16_clk),
    .D(_0223_),
    .Q(\ram[32][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3662_ (.CLK(clknet_leaf_12_clk),
    .D(_0224_),
    .Q(\ram[32][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3663_ (.CLK(clknet_leaf_16_clk),
    .D(_0225_),
    .Q(\ram[32][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3664_ (.CLK(clknet_leaf_14_clk),
    .D(_0226_),
    .Q(\ram[32][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3665_ (.CLK(clknet_leaf_15_clk),
    .D(_0227_),
    .Q(\ram[32][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3666_ (.CLK(clknet_leaf_11_clk),
    .D(_0228_),
    .Q(\ram[33][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3667_ (.CLK(clknet_leaf_17_clk),
    .D(_0229_),
    .Q(\ram[33][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3668_ (.CLK(clknet_leaf_11_clk),
    .D(_0230_),
    .Q(\ram[33][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3669_ (.CLK(clknet_leaf_11_clk),
    .D(_0231_),
    .Q(\ram[33][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3670_ (.CLK(clknet_leaf_11_clk),
    .D(_0232_),
    .Q(\ram[33][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3671_ (.CLK(clknet_leaf_12_clk),
    .D(_0233_),
    .Q(\ram[33][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3672_ (.CLK(clknet_leaf_14_clk),
    .D(_0234_),
    .Q(\ram[33][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3673_ (.CLK(clknet_leaf_15_clk),
    .D(_0235_),
    .Q(\ram[33][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3674_ (.CLK(clknet_leaf_11_clk),
    .D(_0236_),
    .Q(\ram[34][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3675_ (.CLK(clknet_leaf_11_clk),
    .D(_0237_),
    .Q(\ram[34][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3676_ (.CLK(clknet_leaf_11_clk),
    .D(_0238_),
    .Q(\ram[34][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3677_ (.CLK(clknet_leaf_11_clk),
    .D(_0239_),
    .Q(\ram[34][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3678_ (.CLK(clknet_leaf_11_clk),
    .D(_0240_),
    .Q(\ram[34][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3679_ (.CLK(clknet_leaf_12_clk),
    .D(_0241_),
    .Q(\ram[34][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3680_ (.CLK(clknet_leaf_14_clk),
    .D(_0242_),
    .Q(\ram[34][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3681_ (.CLK(clknet_leaf_14_clk),
    .D(_0243_),
    .Q(\ram[34][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3682_ (.CLK(clknet_leaf_11_clk),
    .D(_0244_),
    .Q(\ram[35][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3683_ (.CLK(clknet_leaf_11_clk),
    .D(_0245_),
    .Q(\ram[35][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3684_ (.CLK(clknet_leaf_11_clk),
    .D(_0246_),
    .Q(\ram[35][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3685_ (.CLK(clknet_leaf_11_clk),
    .D(_0247_),
    .Q(\ram[35][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3686_ (.CLK(clknet_leaf_11_clk),
    .D(_0248_),
    .Q(\ram[35][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3687_ (.CLK(clknet_leaf_12_clk),
    .D(_0249_),
    .Q(\ram[35][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3688_ (.CLK(clknet_leaf_13_clk),
    .D(_0250_),
    .Q(\ram[35][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3689_ (.CLK(clknet_leaf_13_clk),
    .D(_0251_),
    .Q(\ram[35][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3690_ (.CLK(clknet_leaf_16_clk),
    .D(_0252_),
    .Q(\ram[36][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3691_ (.CLK(clknet_leaf_17_clk),
    .D(_0253_),
    .Q(\ram[36][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3692_ (.CLK(clknet_leaf_16_clk),
    .D(_0254_),
    .Q(\ram[36][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3693_ (.CLK(clknet_leaf_16_clk),
    .D(_0255_),
    .Q(\ram[36][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3694_ (.CLK(clknet_leaf_16_clk),
    .D(_0256_),
    .Q(\ram[36][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3695_ (.CLK(clknet_leaf_15_clk),
    .D(_0257_),
    .Q(\ram[36][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3696_ (.CLK(clknet_leaf_14_clk),
    .D(_0258_),
    .Q(\ram[36][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3697_ (.CLK(clknet_leaf_15_clk),
    .D(_0259_),
    .Q(\ram[36][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3698_ (.CLK(clknet_leaf_19_clk),
    .D(_0260_),
    .Q(\ram[37][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3699_ (.CLK(clknet_leaf_19_clk),
    .D(_0261_),
    .Q(\ram[37][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3700_ (.CLK(clknet_leaf_18_clk),
    .D(_0262_),
    .Q(\ram[37][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3701_ (.CLK(clknet_leaf_18_clk),
    .D(_0263_),
    .Q(\ram[37][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3702_ (.CLK(clknet_leaf_19_clk),
    .D(_0264_),
    .Q(\ram[37][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3703_ (.CLK(clknet_leaf_21_clk),
    .D(_0265_),
    .Q(\ram[37][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3704_ (.CLK(clknet_leaf_24_clk),
    .D(_0266_),
    .Q(\ram[37][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3705_ (.CLK(clknet_leaf_23_clk),
    .D(_0267_),
    .Q(\ram[37][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3706_ (.CLK(clknet_leaf_17_clk),
    .D(_0268_),
    .Q(\ram[38][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3707_ (.CLK(clknet_leaf_17_clk),
    .D(_0269_),
    .Q(\ram[38][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3708_ (.CLK(clknet_leaf_16_clk),
    .D(_0270_),
    .Q(\ram[38][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3709_ (.CLK(clknet_leaf_18_clk),
    .D(_0271_),
    .Q(\ram[38][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3710_ (.CLK(clknet_leaf_15_clk),
    .D(_0272_),
    .Q(\ram[38][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3711_ (.CLK(clknet_leaf_15_clk),
    .D(_0273_),
    .Q(\ram[38][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3712_ (.CLK(clknet_leaf_25_clk),
    .D(_0274_),
    .Q(\ram[38][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3713_ (.CLK(clknet_leaf_15_clk),
    .D(_0275_),
    .Q(\ram[38][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3714_ (.CLK(clknet_leaf_42_clk),
    .D(_0276_),
    .Q(\ram[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3715_ (.CLK(clknet_leaf_44_clk),
    .D(_0277_),
    .Q(\ram[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3716_ (.CLK(clknet_leaf_41_clk),
    .D(_0278_),
    .Q(\ram[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3717_ (.CLK(clknet_leaf_40_clk),
    .D(_0279_),
    .Q(\ram[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3718_ (.CLK(clknet_leaf_41_clk),
    .D(_0280_),
    .Q(\ram[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3719_ (.CLK(clknet_leaf_41_clk),
    .D(_0281_),
    .Q(\ram[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3720_ (.CLK(clknet_leaf_35_clk),
    .D(_0282_),
    .Q(\ram[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3721_ (.CLK(clknet_leaf_37_clk),
    .D(_0283_),
    .Q(\ram[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3722_ (.CLK(clknet_leaf_17_clk),
    .D(_0284_),
    .Q(\ram[40][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3723_ (.CLK(clknet_leaf_17_clk),
    .D(_0285_),
    .Q(\ram[40][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3724_ (.CLK(clknet_leaf_17_clk),
    .D(_0286_),
    .Q(\ram[40][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3725_ (.CLK(clknet_leaf_17_clk),
    .D(_0287_),
    .Q(\ram[40][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3726_ (.CLK(clknet_leaf_15_clk),
    .D(_0288_),
    .Q(\ram[40][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3727_ (.CLK(clknet_leaf_15_clk),
    .D(_0289_),
    .Q(\ram[40][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3728_ (.CLK(clknet_leaf_24_clk),
    .D(_0290_),
    .Q(\ram[40][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3729_ (.CLK(clknet_leaf_15_clk),
    .D(_0291_),
    .Q(\ram[40][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3730_ (.CLK(clknet_leaf_18_clk),
    .D(_0292_),
    .Q(\ram[41][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3731_ (.CLK(clknet_leaf_17_clk),
    .D(_0293_),
    .Q(\ram[41][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3732_ (.CLK(clknet_leaf_17_clk),
    .D(_0294_),
    .Q(\ram[41][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3733_ (.CLK(clknet_leaf_18_clk),
    .D(_0295_),
    .Q(\ram[41][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3734_ (.CLK(clknet_leaf_18_clk),
    .D(_0296_),
    .Q(\ram[41][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3735_ (.CLK(clknet_leaf_24_clk),
    .D(_0297_),
    .Q(\ram[41][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3736_ (.CLK(clknet_leaf_25_clk),
    .D(_0298_),
    .Q(\ram[41][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3737_ (.CLK(clknet_leaf_24_clk),
    .D(_0299_),
    .Q(\ram[41][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3738_ (.CLK(clknet_leaf_19_clk),
    .D(_0300_),
    .Q(\ram[42][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3739_ (.CLK(clknet_leaf_19_clk),
    .D(_0301_),
    .Q(\ram[42][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3740_ (.CLK(clknet_leaf_19_clk),
    .D(_0302_),
    .Q(\ram[42][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3741_ (.CLK(clknet_leaf_19_clk),
    .D(_0303_),
    .Q(\ram[42][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3742_ (.CLK(clknet_leaf_20_clk),
    .D(_0304_),
    .Q(\ram[42][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3743_ (.CLK(clknet_leaf_21_clk),
    .D(_0305_),
    .Q(\ram[42][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3744_ (.CLK(clknet_leaf_23_clk),
    .D(_0306_),
    .Q(\ram[42][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3745_ (.CLK(clknet_leaf_21_clk),
    .D(_0307_),
    .Q(\ram[42][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3746_ (.CLK(clknet_leaf_19_clk),
    .D(_0308_),
    .Q(\ram[43][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3747_ (.CLK(clknet_leaf_19_clk),
    .D(_0309_),
    .Q(\ram[43][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3748_ (.CLK(clknet_leaf_19_clk),
    .D(_0310_),
    .Q(\ram[43][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3749_ (.CLK(clknet_leaf_19_clk),
    .D(_0311_),
    .Q(\ram[43][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3750_ (.CLK(clknet_leaf_20_clk),
    .D(_0312_),
    .Q(\ram[43][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3751_ (.CLK(clknet_leaf_21_clk),
    .D(_0313_),
    .Q(\ram[43][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3752_ (.CLK(clknet_leaf_21_clk),
    .D(_0314_),
    .Q(\ram[43][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3753_ (.CLK(clknet_leaf_21_clk),
    .D(_0315_),
    .Q(\ram[43][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3754_ (.CLK(clknet_leaf_20_clk),
    .D(_0316_),
    .Q(\ram[44][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3755_ (.CLK(clknet_leaf_20_clk),
    .D(_0317_),
    .Q(\ram[44][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3756_ (.CLK(clknet_leaf_20_clk),
    .D(_0318_),
    .Q(\ram[44][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3757_ (.CLK(clknet_leaf_20_clk),
    .D(_0319_),
    .Q(\ram[44][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3758_ (.CLK(clknet_leaf_20_clk),
    .D(_0320_),
    .Q(\ram[44][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3759_ (.CLK(clknet_leaf_21_clk),
    .D(_0321_),
    .Q(\ram[44][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3760_ (.CLK(clknet_leaf_22_clk),
    .D(_0322_),
    .Q(\ram[44][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3761_ (.CLK(clknet_leaf_22_clk),
    .D(_0323_),
    .Q(\ram[44][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3762_ (.CLK(clknet_leaf_20_clk),
    .D(_0324_),
    .Q(\ram[45][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3763_ (.CLK(clknet_leaf_19_clk),
    .D(_0325_),
    .Q(\ram[45][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3764_ (.CLK(clknet_leaf_20_clk),
    .D(_0326_),
    .Q(\ram[45][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3765_ (.CLK(clknet_leaf_20_clk),
    .D(_0327_),
    .Q(\ram[45][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3766_ (.CLK(clknet_leaf_20_clk),
    .D(_0328_),
    .Q(\ram[45][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3767_ (.CLK(clknet_leaf_21_clk),
    .D(_0329_),
    .Q(\ram[45][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3768_ (.CLK(clknet_leaf_22_clk),
    .D(_0330_),
    .Q(\ram[45][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3769_ (.CLK(clknet_leaf_22_clk),
    .D(_0331_),
    .Q(\ram[45][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3770_ (.CLK(clknet_leaf_20_clk),
    .D(_0332_),
    .Q(\ram[46][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3771_ (.CLK(clknet_leaf_19_clk),
    .D(_0333_),
    .Q(\ram[46][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3772_ (.CLK(clknet_leaf_20_clk),
    .D(_0334_),
    .Q(\ram[46][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3773_ (.CLK(clknet_leaf_20_clk),
    .D(_0335_),
    .Q(\ram[46][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3774_ (.CLK(clknet_leaf_20_clk),
    .D(_0336_),
    .Q(\ram[46][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3775_ (.CLK(clknet_leaf_21_clk),
    .D(_0337_),
    .Q(\ram[46][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3776_ (.CLK(clknet_leaf_22_clk),
    .D(_0338_),
    .Q(\ram[46][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3777_ (.CLK(clknet_leaf_22_clk),
    .D(_0339_),
    .Q(\ram[46][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3778_ (.CLK(clknet_leaf_20_clk),
    .D(_0340_),
    .Q(\ram[47][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3779_ (.CLK(clknet_leaf_19_clk),
    .D(_0341_),
    .Q(\ram[47][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3780_ (.CLK(clknet_leaf_20_clk),
    .D(_0342_),
    .Q(\ram[47][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3781_ (.CLK(clknet_leaf_20_clk),
    .D(_0343_),
    .Q(\ram[47][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3782_ (.CLK(clknet_leaf_20_clk),
    .D(_0344_),
    .Q(\ram[47][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3783_ (.CLK(clknet_leaf_21_clk),
    .D(_0345_),
    .Q(\ram[47][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3784_ (.CLK(clknet_leaf_22_clk),
    .D(_0346_),
    .Q(\ram[47][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3785_ (.CLK(clknet_leaf_22_clk),
    .D(_0347_),
    .Q(\ram[47][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3786_ (.CLK(clknet_leaf_36_clk),
    .D(_0348_),
    .Q(\ram[48][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3787_ (.CLK(clknet_leaf_27_clk),
    .D(_0349_),
    .Q(\ram[48][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3788_ (.CLK(clknet_leaf_36_clk),
    .D(_0350_),
    .Q(\ram[48][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3789_ (.CLK(clknet_leaf_36_clk),
    .D(_0351_),
    .Q(\ram[48][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3790_ (.CLK(clknet_leaf_36_clk),
    .D(_0352_),
    .Q(\ram[48][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3791_ (.CLK(clknet_leaf_27_clk),
    .D(_0353_),
    .Q(\ram[48][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3792_ (.CLK(clknet_leaf_25_clk),
    .D(_0354_),
    .Q(\ram[48][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3793_ (.CLK(clknet_leaf_25_clk),
    .D(_0355_),
    .Q(\ram[48][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3794_ (.CLK(clknet_leaf_40_clk),
    .D(_0356_),
    .Q(\ram[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3795_ (.CLK(clknet_leaf_39_clk),
    .D(_0357_),
    .Q(\ram[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3796_ (.CLK(clknet_leaf_35_clk),
    .D(_0358_),
    .Q(\ram[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3797_ (.CLK(clknet_leaf_40_clk),
    .D(_0359_),
    .Q(\ram[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3798_ (.CLK(clknet_leaf_40_clk),
    .D(_0360_),
    .Q(\ram[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3799_ (.CLK(clknet_leaf_35_clk),
    .D(_0361_),
    .Q(\ram[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3800_ (.CLK(clknet_leaf_37_clk),
    .D(_0362_),
    .Q(\ram[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3801_ (.CLK(clknet_leaf_37_clk),
    .D(_0363_),
    .Q(\ram[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3802_ (.CLK(clknet_leaf_23_clk),
    .D(_0364_),
    .Q(\ram[50][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3803_ (.CLK(clknet_leaf_23_clk),
    .D(_0365_),
    .Q(\ram[50][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3804_ (.CLK(clknet_leaf_23_clk),
    .D(_0366_),
    .Q(\ram[50][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3805_ (.CLK(clknet_leaf_23_clk),
    .D(_0367_),
    .Q(\ram[50][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3806_ (.CLK(clknet_leaf_23_clk),
    .D(_0368_),
    .Q(\ram[50][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3807_ (.CLK(clknet_leaf_23_clk),
    .D(_0369_),
    .Q(\ram[50][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3808_ (.CLK(clknet_leaf_23_clk),
    .D(_0370_),
    .Q(\ram[50][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3809_ (.CLK(clknet_leaf_23_clk),
    .D(_0371_),
    .Q(\ram[50][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3810_ (.CLK(clknet_leaf_28_clk),
    .D(_0372_),
    .Q(\ram[51][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3811_ (.CLK(clknet_leaf_28_clk),
    .D(_0373_),
    .Q(\ram[51][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3812_ (.CLK(clknet_leaf_30_clk),
    .D(_0374_),
    .Q(\ram[51][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3813_ (.CLK(clknet_leaf_28_clk),
    .D(_0375_),
    .Q(\ram[51][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3814_ (.CLK(clknet_leaf_30_clk),
    .D(_0376_),
    .Q(\ram[51][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3815_ (.CLK(clknet_leaf_28_clk),
    .D(_0377_),
    .Q(\ram[51][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3816_ (.CLK(clknet_leaf_23_clk),
    .D(_0378_),
    .Q(\ram[51][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3817_ (.CLK(clknet_leaf_23_clk),
    .D(_0379_),
    .Q(\ram[51][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3818_ (.CLK(clknet_leaf_29_clk),
    .D(_0380_),
    .Q(\ram[52][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3819_ (.CLK(clknet_leaf_29_clk),
    .D(_0381_),
    .Q(\ram[52][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3820_ (.CLK(clknet_leaf_30_clk),
    .D(_0382_),
    .Q(\ram[52][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3821_ (.CLK(clknet_leaf_30_clk),
    .D(_0383_),
    .Q(\ram[52][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3822_ (.CLK(clknet_leaf_31_clk),
    .D(_0384_),
    .Q(\ram[52][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3823_ (.CLK(clknet_leaf_30_clk),
    .D(_0385_),
    .Q(\ram[52][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3824_ (.CLK(clknet_leaf_23_clk),
    .D(_0386_),
    .Q(\ram[52][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3825_ (.CLK(clknet_leaf_22_clk),
    .D(_0387_),
    .Q(\ram[52][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3826_ (.CLK(clknet_leaf_29_clk),
    .D(_0388_),
    .Q(\ram[53][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3827_ (.CLK(clknet_leaf_29_clk),
    .D(_0389_),
    .Q(\ram[53][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3828_ (.CLK(clknet_leaf_31_clk),
    .D(_0390_),
    .Q(\ram[53][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3829_ (.CLK(clknet_leaf_29_clk),
    .D(_0391_),
    .Q(\ram[53][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3830_ (.CLK(clknet_leaf_31_clk),
    .D(_0392_),
    .Q(\ram[53][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3831_ (.CLK(clknet_leaf_30_clk),
    .D(_0393_),
    .Q(\ram[53][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3832_ (.CLK(clknet_leaf_29_clk),
    .D(_0394_),
    .Q(\ram[53][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3833_ (.CLK(clknet_leaf_29_clk),
    .D(_0395_),
    .Q(\ram[53][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3834_ (.CLK(clknet_leaf_29_clk),
    .D(_0396_),
    .Q(\ram[54][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3835_ (.CLK(clknet_leaf_28_clk),
    .D(_0397_),
    .Q(\ram[54][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3836_ (.CLK(clknet_leaf_31_clk),
    .D(_0398_),
    .Q(\ram[54][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3837_ (.CLK(clknet_leaf_30_clk),
    .D(_0399_),
    .Q(\ram[54][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3838_ (.CLK(clknet_leaf_31_clk),
    .D(_0400_),
    .Q(\ram[54][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3839_ (.CLK(clknet_leaf_30_clk),
    .D(_0401_),
    .Q(\ram[54][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3840_ (.CLK(clknet_leaf_29_clk),
    .D(_0402_),
    .Q(\ram[54][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3841_ (.CLK(clknet_leaf_22_clk),
    .D(_0403_),
    .Q(\ram[54][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3842_ (.CLK(clknet_leaf_29_clk),
    .D(_0404_),
    .Q(\ram[55][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3843_ (.CLK(clknet_leaf_29_clk),
    .D(_0405_),
    .Q(\ram[55][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3844_ (.CLK(clknet_leaf_31_clk),
    .D(_0406_),
    .Q(\ram[55][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3845_ (.CLK(clknet_leaf_30_clk),
    .D(_0407_),
    .Q(\ram[55][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3846_ (.CLK(clknet_leaf_31_clk),
    .D(_0408_),
    .Q(\ram[55][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3847_ (.CLK(clknet_leaf_30_clk),
    .D(_0409_),
    .Q(\ram[55][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3848_ (.CLK(clknet_leaf_29_clk),
    .D(_0410_),
    .Q(\ram[55][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3849_ (.CLK(clknet_leaf_22_clk),
    .D(_0411_),
    .Q(\ram[55][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3850_ (.CLK(clknet_leaf_36_clk),
    .D(_0412_),
    .Q(\ram[56][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3851_ (.CLK(clknet_leaf_36_clk),
    .D(_0413_),
    .Q(\ram[56][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3852_ (.CLK(clknet_leaf_33_clk),
    .D(_0414_),
    .Q(\ram[56][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3853_ (.CLK(clknet_leaf_34_clk),
    .D(_0415_),
    .Q(\ram[56][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3854_ (.CLK(clknet_leaf_34_clk),
    .D(_0416_),
    .Q(\ram[56][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3855_ (.CLK(clknet_leaf_33_clk),
    .D(_0417_),
    .Q(\ram[56][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3856_ (.CLK(clknet_leaf_27_clk),
    .D(_0418_),
    .Q(\ram[56][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3857_ (.CLK(clknet_leaf_27_clk),
    .D(_0419_),
    .Q(\ram[56][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3858_ (.CLK(clknet_leaf_36_clk),
    .D(_0420_),
    .Q(\ram[57][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3859_ (.CLK(clknet_leaf_36_clk),
    .D(_0421_),
    .Q(\ram[57][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3860_ (.CLK(clknet_leaf_35_clk),
    .D(_0422_),
    .Q(\ram[57][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3861_ (.CLK(clknet_leaf_34_clk),
    .D(_0423_),
    .Q(\ram[57][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3862_ (.CLK(clknet_leaf_34_clk),
    .D(_0424_),
    .Q(\ram[57][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3863_ (.CLK(clknet_leaf_33_clk),
    .D(_0425_),
    .Q(\ram[57][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3864_ (.CLK(clknet_leaf_26_clk),
    .D(_0426_),
    .Q(\ram[57][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3865_ (.CLK(clknet_leaf_27_clk),
    .D(_0427_),
    .Q(\ram[57][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3866_ (.CLK(clknet_leaf_35_clk),
    .D(_0428_),
    .Q(\ram[58][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3867_ (.CLK(clknet_leaf_36_clk),
    .D(_0429_),
    .Q(\ram[58][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3868_ (.CLK(clknet_leaf_35_clk),
    .D(_0430_),
    .Q(\ram[58][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3869_ (.CLK(clknet_leaf_34_clk),
    .D(_0431_),
    .Q(\ram[58][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3870_ (.CLK(clknet_leaf_34_clk),
    .D(_0432_),
    .Q(\ram[58][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3871_ (.CLK(clknet_leaf_33_clk),
    .D(_0433_),
    .Q(\ram[58][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3872_ (.CLK(clknet_leaf_26_clk),
    .D(_0434_),
    .Q(\ram[58][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3873_ (.CLK(clknet_leaf_27_clk),
    .D(_0435_),
    .Q(\ram[58][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3874_ (.CLK(clknet_leaf_40_clk),
    .D(_0436_),
    .Q(\ram[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3875_ (.CLK(clknet_leaf_39_clk),
    .D(_0437_),
    .Q(\ram[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3876_ (.CLK(clknet_leaf_35_clk),
    .D(_0438_),
    .Q(\ram[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3877_ (.CLK(clknet_leaf_40_clk),
    .D(_0439_),
    .Q(\ram[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3878_ (.CLK(clknet_leaf_35_clk),
    .D(_0440_),
    .Q(\ram[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3879_ (.CLK(clknet_leaf_35_clk),
    .D(_0441_),
    .Q(\ram[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3880_ (.CLK(clknet_leaf_36_clk),
    .D(_0442_),
    .Q(\ram[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3881_ (.CLK(clknet_leaf_37_clk),
    .D(_0443_),
    .Q(\ram[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3882_ (.CLK(clknet_leaf_30_clk),
    .D(_0444_),
    .Q(\ram[60][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3883_ (.CLK(clknet_leaf_30_clk),
    .D(_0445_),
    .Q(\ram[60][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3884_ (.CLK(clknet_leaf_31_clk),
    .D(_0446_),
    .Q(\ram[60][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3885_ (.CLK(clknet_leaf_32_clk),
    .D(_0447_),
    .Q(\ram[60][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3886_ (.CLK(clknet_leaf_32_clk),
    .D(_0448_),
    .Q(\ram[60][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3887_ (.CLK(clknet_leaf_32_clk),
    .D(_0449_),
    .Q(\ram[60][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3888_ (.CLK(clknet_leaf_28_clk),
    .D(_0450_),
    .Q(\ram[60][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3889_ (.CLK(clknet_leaf_28_clk),
    .D(_0451_),
    .Q(\ram[60][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3890_ (.CLK(clknet_leaf_30_clk),
    .D(_0452_),
    .Q(\ram[61][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3891_ (.CLK(clknet_leaf_30_clk),
    .D(_0453_),
    .Q(\ram[61][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3892_ (.CLK(clknet_leaf_32_clk),
    .D(_0454_),
    .Q(\ram[61][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3893_ (.CLK(clknet_leaf_31_clk),
    .D(_0455_),
    .Q(\ram[61][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3894_ (.CLK(clknet_leaf_32_clk),
    .D(_0456_),
    .Q(\ram[61][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3895_ (.CLK(clknet_leaf_30_clk),
    .D(_0457_),
    .Q(\ram[61][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3896_ (.CLK(clknet_leaf_28_clk),
    .D(_0458_),
    .Q(\ram[61][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3897_ (.CLK(clknet_leaf_28_clk),
    .D(_0459_),
    .Q(\ram[61][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3898_ (.CLK(clknet_leaf_32_clk),
    .D(_0460_),
    .Q(\ram[62][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3899_ (.CLK(clknet_leaf_33_clk),
    .D(_0461_),
    .Q(\ram[62][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3900_ (.CLK(clknet_leaf_32_clk),
    .D(_0462_),
    .Q(\ram[62][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3901_ (.CLK(clknet_leaf_32_clk),
    .D(_0463_),
    .Q(\ram[62][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3902_ (.CLK(clknet_leaf_32_clk),
    .D(_0464_),
    .Q(\ram[62][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3903_ (.CLK(clknet_leaf_32_clk),
    .D(_0465_),
    .Q(\ram[62][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3904_ (.CLK(clknet_leaf_28_clk),
    .D(_0466_),
    .Q(\ram[62][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3905_ (.CLK(clknet_leaf_28_clk),
    .D(_0467_),
    .Q(\ram[62][7] ));
 sky130_fd_sc_hd__dfxtp_2 _3906_ (.CLK(clknet_leaf_37_clk),
    .D(_0006_),
    .Q(_0000_));
 sky130_fd_sc_hd__dfxtp_1 _3907_ (.CLK(clknet_leaf_26_clk),
    .D(_0007_),
    .Q(_0001_));
 sky130_fd_sc_hd__dfxtp_1 _3908_ (.CLK(clknet_leaf_26_clk),
    .D(_0008_),
    .Q(_0002_));
 sky130_fd_sc_hd__dfxtp_2 _3909_ (.CLK(clknet_leaf_14_clk),
    .D(_0009_),
    .Q(_0003_));
 sky130_fd_sc_hd__dfxtp_4 _3910_ (.CLK(clknet_leaf_14_clk),
    .D(_0010_),
    .Q(_0004_));
 sky130_fd_sc_hd__dfxtp_2 _3911_ (.CLK(clknet_leaf_25_clk),
    .D(_0011_),
    .Q(_0005_));
 sky130_fd_sc_hd__dfxtp_1 _3912_ (.CLK(clknet_leaf_4_clk),
    .D(_0468_),
    .Q(\ram[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3913_ (.CLK(clknet_leaf_10_clk),
    .D(_0469_),
    .Q(\ram[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3914_ (.CLK(clknet_leaf_12_clk),
    .D(_0470_),
    .Q(\ram[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3915_ (.CLK(clknet_leaf_12_clk),
    .D(_0471_),
    .Q(\ram[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3916_ (.CLK(clknet_leaf_12_clk),
    .D(_0472_),
    .Q(\ram[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3917_ (.CLK(clknet_leaf_4_clk),
    .D(_0473_),
    .Q(\ram[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3918_ (.CLK(clknet_leaf_14_clk),
    .D(_0474_),
    .Q(\ram[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3919_ (.CLK(clknet_leaf_13_clk),
    .D(_0475_),
    .Q(\ram[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3920_ (.CLK(clknet_leaf_39_clk),
    .D(_0476_),
    .Q(\ram[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3921_ (.CLK(clknet_leaf_38_clk),
    .D(_0477_),
    .Q(\ram[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3922_ (.CLK(clknet_leaf_41_clk),
    .D(_0478_),
    .Q(\ram[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3923_ (.CLK(clknet_leaf_40_clk),
    .D(_0479_),
    .Q(\ram[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3924_ (.CLK(clknet_leaf_41_clk),
    .D(_0480_),
    .Q(\ram[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3925_ (.CLK(clknet_leaf_39_clk),
    .D(_0481_),
    .Q(\ram[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3926_ (.CLK(clknet_leaf_37_clk),
    .D(_0482_),
    .Q(\ram[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3927_ (.CLK(clknet_leaf_37_clk),
    .D(_0483_),
    .Q(\ram[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3928_ (.CLK(clknet_leaf_33_clk),
    .D(_0484_),
    .Q(\ram[63][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3929_ (.CLK(clknet_leaf_36_clk),
    .D(_0485_),
    .Q(\ram[63][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3930_ (.CLK(clknet_leaf_33_clk),
    .D(_0486_),
    .Q(\ram[63][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3931_ (.CLK(clknet_leaf_32_clk),
    .D(_0487_),
    .Q(\ram[63][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3932_ (.CLK(clknet_leaf_34_clk),
    .D(_0488_),
    .Q(\ram[63][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3933_ (.CLK(clknet_leaf_33_clk),
    .D(_0489_),
    .Q(\ram[63][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3934_ (.CLK(clknet_leaf_28_clk),
    .D(_0490_),
    .Q(\ram[63][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3935_ (.CLK(clknet_leaf_28_clk),
    .D(_0491_),
    .Q(\ram[63][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3936_ (.CLK(clknet_leaf_35_clk),
    .D(_0492_),
    .Q(\ram[59][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3937_ (.CLK(clknet_leaf_36_clk),
    .D(_0493_),
    .Q(\ram[59][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3938_ (.CLK(clknet_leaf_35_clk),
    .D(_0494_),
    .Q(\ram[59][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3939_ (.CLK(clknet_leaf_34_clk),
    .D(_0495_),
    .Q(\ram[59][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3940_ (.CLK(clknet_leaf_34_clk),
    .D(_0496_),
    .Q(\ram[59][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3941_ (.CLK(clknet_leaf_36_clk),
    .D(_0497_),
    .Q(\ram[59][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3942_ (.CLK(clknet_leaf_26_clk),
    .D(_0498_),
    .Q(\ram[59][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3943_ (.CLK(clknet_leaf_27_clk),
    .D(_0499_),
    .Q(\ram[59][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3944_ (.CLK(clknet_leaf_27_clk),
    .D(_0500_),
    .Q(\ram[49][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3945_ (.CLK(clknet_leaf_27_clk),
    .D(_0501_),
    .Q(\ram[49][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3946_ (.CLK(clknet_leaf_36_clk),
    .D(_0502_),
    .Q(\ram[49][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3947_ (.CLK(clknet_leaf_30_clk),
    .D(_0503_),
    .Q(\ram[49][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3948_ (.CLK(clknet_leaf_27_clk),
    .D(_0504_),
    .Q(\ram[49][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3949_ (.CLK(clknet_leaf_27_clk),
    .D(_0505_),
    .Q(\ram[49][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3950_ (.CLK(clknet_leaf_23_clk),
    .D(_0506_),
    .Q(\ram[49][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3951_ (.CLK(clknet_leaf_25_clk),
    .D(_0507_),
    .Q(\ram[49][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3952_ (.CLK(clknet_leaf_43_clk),
    .D(_0508_),
    .Q(\ram[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3953_ (.CLK(clknet_leaf_44_clk),
    .D(_0509_),
    .Q(\ram[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3954_ (.CLK(clknet_leaf_43_clk),
    .D(_0510_),
    .Q(\ram[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3955_ (.CLK(clknet_leaf_42_clk),
    .D(_0511_),
    .Q(\ram[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3956_ (.CLK(clknet_leaf_43_clk),
    .D(_0512_),
    .Q(\ram[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3957_ (.CLK(clknet_leaf_43_clk),
    .D(_0513_),
    .Q(\ram[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3958_ (.CLK(clknet_leaf_39_clk),
    .D(_0514_),
    .Q(\ram[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3959_ (.CLK(clknet_leaf_38_clk),
    .D(_0515_),
    .Q(\ram[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3960_ (.CLK(clknet_leaf_16_clk),
    .D(_0516_),
    .Q(\ram[39][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3961_ (.CLK(clknet_leaf_16_clk),
    .D(_0517_),
    .Q(\ram[39][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3962_ (.CLK(clknet_leaf_16_clk),
    .D(_0518_),
    .Q(\ram[39][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3963_ (.CLK(clknet_leaf_15_clk),
    .D(_0519_),
    .Q(\ram[39][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3964_ (.CLK(clknet_leaf_16_clk),
    .D(_0520_),
    .Q(\ram[39][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3965_ (.CLK(clknet_leaf_15_clk),
    .D(_0521_),
    .Q(\ram[39][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3966_ (.CLK(clknet_leaf_25_clk),
    .D(_0522_),
    .Q(\ram[39][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3967_ (.CLK(clknet_leaf_15_clk),
    .D(_0523_),
    .Q(\ram[39][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3968_ (.CLK(clknet_leaf_37_clk),
    .D(_0524_),
    .Q(\addr_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3969_ (.CLK(clknet_leaf_37_clk),
    .D(_0525_),
    .Q(\addr_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3970_ (.CLK(clknet_leaf_37_clk),
    .D(_0526_),
    .Q(\addr_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3971_ (.CLK(clknet_leaf_14_clk),
    .D(_0527_),
    .Q(\addr_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3972_ (.CLK(clknet_leaf_14_clk),
    .D(_0528_),
    .Q(\addr_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3973_ (.CLK(clknet_leaf_26_clk),
    .D(_0529_),
    .Q(\addr_reg[5] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_10_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_11_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_12_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_13_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_21_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_22_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_23_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_24_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_25_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_26_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_27_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_28_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_29_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_30_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_31_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_32_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_33_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_34_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_35_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_36_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_37_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_38_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_39_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_3_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_40_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_41_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_42_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_43_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_44_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_4_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_5_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_6_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_8_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\addr_reg[5] ),
    .X(net24));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\ram[39][6] ),
    .X(net33));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\ram[22][2] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\ram[63][2] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\ram[40][0] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\ram[32][5] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\ram[22][7] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\ram[28][7] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\ram[15][4] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\ram[20][3] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\ram[58][4] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\ram[36][6] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\ram[16][6] ),
    .X(net34));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\ram[5][0] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\ram[29][2] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\ram[3][2] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\ram[1][2] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\ram[0][0] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\ram[17][2] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\ram[46][5] ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\ram[26][1] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\ram[17][0] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\ram[38][2] ),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\ram[57][6] ),
    .X(net35));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\ram[30][2] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\ram[55][2] ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\ram[24][0] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\ram[0][2] ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\ram[63][5] ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\ram[1][4] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\ram[26][3] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\ram[6][4] ),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\ram[4][2] ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\ram[40][7] ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\ram[25][7] ),
    .X(net36));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\ram[26][4] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\ram[5][1] ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\ram[17][4] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\ram[4][5] ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\ram[44][6] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\ram[1][6] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\ram[6][5] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\ram[7][1] ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\ram[14][6] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\ram[32][6] ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\ram[15][1] ),
    .X(net37));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\ram[2][6] ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\ram[3][6] ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\ram[22][4] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\ram[24][5] ),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\ram[31][2] ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\ram[58][3] ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\ram[20][7] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\ram[8][0] ),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\ram[6][3] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\ram[31][4] ),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\ram[48][7] ),
    .X(net38));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\ram[57][5] ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\ram[24][4] ),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\ram[6][0] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\ram[17][1] ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\ram[0][1] ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\ram[10][7] ),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\ram[32][0] ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\ram[47][5] ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\ram[19][3] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\ram[5][5] ),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\ram[24][6] ),
    .X(net39));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\ram[36][0] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\ram[26][0] ),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\ram[44][7] ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\ram[16][5] ),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\ram[33][3] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\ram[59][0] ),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\ram[43][7] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\ram[23][1] ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\ram[39][4] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\ram[3][5] ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\ram[13][2] ),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\ram[59][4] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\ram[54][0] ),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\ram[9][4] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\ram[40][3] ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\addr_reg[3] ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\ram[26][5] ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\ram[21][4] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\ram[42][5] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\ram[36][5] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\ram[33][6] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\ram[18][7] ),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\ram[16][0] ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\ram[6][2] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\ram[7][0] ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\ram[11][7] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\ram[40][5] ),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\ram[6][7] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\ram[29][1] ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\ram[52][4] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\ram[22][3] ),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\ram[14][1] ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\ram[12][1] ),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\ram[36][7] ),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\ram[3][3] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\ram[25][6] ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\ram[21][0] ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\ram[16][4] ),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\ram[2][0] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\ram[29][3] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\ram[3][7] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\ram[15][7] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\ram[1][1] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\ram[40][6] ),
    .X(net25));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\ram[16][7] ),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\ram[53][4] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\ram[12][6] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\ram[53][0] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\ram[26][7] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\ram[5][2] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\ram[57][4] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\ram[54][4] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\ram[14][4] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\ram[9][2] ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\ram[62][0] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\ram[6][1] ),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\ram[62][3] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\ram[62][5] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\ram[62][4] ),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\ram[8][4] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\ram[0][7] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\ram[15][0] ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\ram[33][7] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\ram[57][2] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\ram[13][0] ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\ram[10][6] ),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\ram[38][6] ),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\ram[9][6] ),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\ram[24][1] ),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\ram[35][5] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\ram[4][4] ),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\ram[47][7] ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\ram[22][5] ),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\ram[32][1] ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\ram[58][2] ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\ram[13][7] ),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\ram[43][6] ),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\ram[49][7] ),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\ram[7][5] ),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\ram[52][1] ),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\ram[61][6] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\ram[28][1] ),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\ram[3][4] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\ram[4][0] ),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\ram[22][1] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\ram[26][6] ),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\ram[26][2] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\ram[12][0] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\ram[41][0] ),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\ram[0][4] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\ram[9][7] ),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\ram[30][4] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\ram[30][0] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\ram[4][7] ),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\ram[30][7] ),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\ram[54][1] ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\ram[34][1] ),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\ram[37][5] ),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\ram[48][4] ),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\ram[37][6] ),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\ram[42][2] ),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\ram[33][0] ),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\ram[0][5] ),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\ram[16][1] ),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\ram[10][1] ),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\ram[58][7] ),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\ram[4][6] ),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\ram[31][7] ),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\ram[19][4] ),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\addr_reg[4] ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\ram[20][2] ),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\ram[5][4] ),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\ram[34][2] ),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\ram[30][3] ),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\ram[39][3] ),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\ram[23][6] ),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\ram[13][4] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\ram[7][3] ),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\ram[59][2] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\ram[38][4] ),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\ram[31][1] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\ram[23][7] ),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\ram[1][3] ),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\ram[54][7] ),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\ram[32][3] ),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\ram[19][2] ),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\ram[10][2] ),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\ram[5][3] ),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\ram[40][2] ),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\ram[60][3] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\ram[24][7] ),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\ram[55][1] ),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\ram[8][5] ),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\ram[11][5] ),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\ram[41][2] ),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\ram[21][2] ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\ram[59][3] ),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\ram[36][2] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\ram[40][4] ),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\ram[10][4] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\ram[39][5] ),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\ram[20][5] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\ram[7][7] ),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\ram[8][3] ),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\ram[10][3] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\ram[60][5] ),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\ram[54][6] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\ram[38][0] ),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\ram[51][0] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\ram[18][0] ),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\ram[15][5] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\ram[46][7] ),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\ram[47][1] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\ram[8][7] ),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\ram[41][3] ),
    .X(net26));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\ram[62][1] ),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\ram[48][3] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\ram[43][5] ),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\ram[56][0] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\ram[20][6] ),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\ram[7][6] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\ram[40][1] ),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\ram[22][6] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\ram[33][4] ),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\ram[7][4] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\ram[39][7] ),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\ram[13][1] ),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\ram[42][6] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\ram[57][7] ),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\ram[25][1] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\ram[18][2] ),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\ram[30][6] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\ram[20][1] ),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\ram[51][1] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\ram[41][1] ),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\ram[6][6] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\ram[59][7] ),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\ram[33][5] ),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\ram[13][6] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\ram[39][2] ),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\ram[31][3] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\ram[23][5] ),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\ram[25][5] ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\ram[8][6] ),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\ram[33][2] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\ram[4][3] ),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\ram[21][5] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\ram[34][4] ),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\ram[34][5] ),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\ram[2][4] ),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\ram[42][0] ),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\ram[31][0] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\ram[51][5] ),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(\ram[27][1] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\ram[52][6] ),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\ram[43][3] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\ram[2][5] ),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\ram[53][1] ),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\ram[49][5] ),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\ram[59][6] ),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\ram[7][2] ),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\ram[63][4] ),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\ram[25][2] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\ram[63][6] ),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\ram[56][6] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\ram[45][7] ),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\ram[38][5] ),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\ram[1][7] ),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\ram[34][3] ),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\ram[55][7] ),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\ram[38][3] ),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\ram[18][4] ),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\ram[19][1] ),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(\ram[13][5] ),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\ram[25][0] ),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\ram[31][6] ),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\ram[2][7] ),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\ram[60][7] ),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\ram[15][3] ),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\ram[24][3] ),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\ram[29][7] ),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\ram[34][7] ),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\ram[46][1] ),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\ram[12][7] ),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\addr_reg[1] ),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\ram[12][5] ),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\ram[12][4] ),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\ram[39][1] ),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\ram[38][7] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\ram[8][2] ),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\ram[27][7] ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\ram[10][0] ),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\ram[15][2] ),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\ram[30][5] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\ram[17][3] ),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\ram[42][1] ),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\ram[63][7] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\ram[59][1] ),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\ram[53][3] ),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\ram[19][6] ),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\ram[49][1] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\ram[39][0] ),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\ram[46][6] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\ram[48][6] ),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\ram[60][6] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\ram[29][6] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\ram[55][0] ),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\ram[48][0] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\ram[29][5] ),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\ram[56][1] ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\ram[28][5] ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\ram[18][1] ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\ram[62][6] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\ram[3][1] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\ram[23][0] ),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\ram[59][5] ),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\ram[53][5] ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\ram[51][3] ),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\ram[49][4] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\ram[55][5] ),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\ram[62][2] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\ram[14][0] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\ram[5][7] ),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\ram[14][7] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\ram[48][2] ),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\ram[41][5] ),
    .X(net27));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\ram[45][5] ),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(\ram[58][0] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\ram[61][2] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\ram[18][5] ),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\ram[25][3] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\ram[27][5] ),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\ram[45][4] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\ram[52][7] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\ram[14][3] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(\ram[54][5] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\ram[54][3] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\ram[16][2] ),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(\ram[34][0] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\ram[32][7] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\ram[11][6] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\ram[5][6] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\ram[14][5] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\ram[62][7] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\ram[61][4] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\ram[43][1] ),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\ram[19][0] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\ram[55][3] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\ram[0][3] ),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(\ram[31][5] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\ram[46][2] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(\ram[35][6] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\ram[43][2] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(\ram[49][0] ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\ram[30][1] ),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(\ram[27][6] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\ram[52][0] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(\ram[60][0] ),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\ram[36][3] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\ram[28][3] ),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\ram[38][1] ),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\ram[52][5] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(\ram[61][7] ),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\ram[42][3] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\ram[13][3] ),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\ram[63][3] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\ram[61][3] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\ram[50][7] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\ram[53][6] ),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\ram[12][3] ),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\ram[23][2] ),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\addr_reg[0] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\ram[21][1] ),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\ram[53][7] ),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\ram[27][0] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(\ram[57][1] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\ram[25][4] ),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\ram[42][4] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\ram[45][1] ),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(\ram[44][1] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\ram[35][7] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\ram[56][3] ),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\ram[11][1] ),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\ram[8][1] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\ram[44][0] ),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\addr_reg[2] ),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\ram[37][4] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\ram[60][1] ),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\ram[57][0] ),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\ram[58][1] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\ram[45][3] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\ram[44][3] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\ram[55][4] ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\ram[49][6] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\ram[29][0] ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\ram[46][4] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\ram[27][3] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\ram[27][4] ),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\ram[0][6] ),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\ram[18][3] ),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\ram[11][3] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\ram[52][3] ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\ram[60][4] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\ram[12][2] ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\ram[50][6] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\ram[63][1] ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\ram[32][2] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\ram[49][3] ),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\ram[55][6] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\ram[27][2] ),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\ram[51][6] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\ram[37][7] ),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\ram[45][2] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\ram[35][4] ),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\ram[54][2] ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\ram[52][2] ),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\ram[9][1] ),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\ram[46][0] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\ram[35][3] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\ram[35][0] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\ram[43][4] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\ram[47][4] ),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\ram[47][2] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\ram[51][4] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\ram[45][6] ),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\ram[17][6] ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\ram[24][2] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\ram[46][3] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\ram[61][5] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\ram[47][0] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\ram[37][1] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\ram[45][0] ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\ram[44][4] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\ram[43][0] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\ram[51][2] ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\ram[11][0] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\ram[58][6] ),
    .X(net28));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\ram[56][4] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(\ram[44][2] ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\ram[51][7] ),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(\ram[17][5] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\ram[47][3] ),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(\ram[19][5] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\ram[11][2] ),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\ram[49][2] ),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\ram[11][4] ),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\ram[61][0] ),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\ram[4][1] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\ram[28][4] ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\ram[63][0] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\ram[3][0] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\ram[42][7] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\ram[58][5] ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\ram[57][3] ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\ram[34][6] ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\ram[1][5] ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\ram[1][0] ),
    .X(net29));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\ram[41][4] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\ram[20][4] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\ram[53][2] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\ram[56][5] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\ram[48][5] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\ram[20][0] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\ram[9][5] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\ram[17][7] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\ram[28][2] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\ram[44][5] ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\ram[56][2] ),
    .X(net30));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\ram[36][4] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\ram[10][5] ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\ram[37][3] ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\ram[18][6] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\ram[32][4] ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\ram[19][7] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\ram[41][6] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\ram[23][3] ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\ram[21][7] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\ram[28][6] ),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\ram[15][6] ),
    .X(net31));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\ram[60][2] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\ram[37][2] ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\ram[48][1] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\ram[21][3] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\ram[9][3] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\ram[56][7] ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\ram[14][2] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\ram[16][3] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\ram[9][0] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\ram[36][1] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\ram[41][7] ),
    .X(net32));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\ram[23][4] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\ram[2][3] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\ram[21][6] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\ram[33][1] ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\ram[2][2] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\ram[28][0] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\ram[29][4] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\ram[2][1] ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\ram[22][0] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\ram[47][6] ),
    .X(net122));
 sky130_fd_sc_hd__buf_1 input1 (.A(addr[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input10 (.A(data[3]),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input11 (.A(data[4]),
    .X(net11));
 sky130_fd_sc_hd__buf_4 input12 (.A(data[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(data[6]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(data[7]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input15 (.A(we),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input2 (.A(addr[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(addr[2]),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(addr[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(addr[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(addr[5]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(data[0]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input8 (.A(data[1]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(data[2]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 output16 (.A(net16),
    .X(q[0]));
 sky130_fd_sc_hd__clkbuf_4 output17 (.A(net17),
    .X(q[1]));
 sky130_fd_sc_hd__clkbuf_4 output18 (.A(net18),
    .X(q[2]));
 sky130_fd_sc_hd__clkbuf_4 output19 (.A(net19),
    .X(q[3]));
 sky130_fd_sc_hd__clkbuf_4 output20 (.A(net20),
    .X(q[4]));
 sky130_fd_sc_hd__clkbuf_4 output21 (.A(net21),
    .X(q[5]));
 sky130_fd_sc_hd__clkbuf_4 output22 (.A(net22),
    .X(q[6]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(q[7]));
endmodule

